��z     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�M �estimator_params�(�	criterion��	max_depth��min_samples_split��min_samples_leaf��min_weight_fraction_leaf��max_features��max_leaf_nodes��min_impurity_decrease��random_state��	ccp_alpha�t��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�Nh�entropy�hKhKhKhG        h�auto�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h6�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C`                                                                	       
              �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hh.hhhKhKhKhG        h�sqrt�hNhJ/�LjhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��h?�f8�����R�(KhCNNNJ����J����K t�b�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGh3�scalar���h?�i8�����R�(KhCNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hK�
node_count�K�nodes�h5h8K ��h:��R�(KK��h?�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hyh\K ��hzh\K��h{h\K��h|h?�f8�����R�(KhCNNNJ����J����K t�bK��h}h�K ��h~h\K(��hh�K0��uK8KKt�b�B�                             �?�?�T@�	           ��@       	                   �5@ԭ�3k@           |�@                           �?y"���@�           �@                            @��eP0@�             m@������������������������       ��@�'@V            �_@������������������������       ���ɍZ@D            �Z@                           @ߴS�@G           �@������������������������       �R9�+x@�            @j@������������������������       �б{Hh @�            �r@
                           �?��z��5@%           �{@                           �?����:�@�            `l@������������������������       �1��\@F            �Y@������������������������       �ק9��@I             _@                            �?�<LK�@�             k@������������������������       �>*�F�@             �E@������������������������       ��Y4��d@v            �e@                          �4@k�R��A@�           T�@                          �1@J�]�
@�           T�@                           @H���Q=@�            Pw@������������������������       �k��/�@s             g@������������������������       �Ě/�/��?x            �g@                           @�4�|��@�            �@������������������������       �����@H           p�@������������������������       �W�Tf�@�             q@                           @����]	@�           T�@                          �9@�N?�/H
@c           ��@������������������������       ��7fJ��	@l           ��@������������������������       ����6
@�            �w@                          �8@W_E�jZ@e           �@������������������������       ���^��<@�            �w@������������������������       �����@�            �l@�t�b�values�h5h8K ��h:��R�(KKKK��h��B�        4@     �s@     ��@      A@      L@     `{@     @W@     ��@     @i@      �@     �v@      >@             �W@     �c@       @      @     �[@      $@     `z@      A@     �p@     @S@      @              F@     �V@       @             �K@      @     pt@      7@     �c@     �@@      �?              4@      ?@       @              8@      �?      T@      .@      F@      .@      �?              &@      *@       @              *@      �?     �B@      &@      <@      "@      �?              "@      2@                      &@             �E@      @      0@      @                      8@     �M@                      ?@      @     �n@       @     �\@      2@                      ,@      ;@                      0@      @     �U@             �M@      @                      $@      @@                      .@              d@       @      L@      ,@                      I@     @Q@              @      L@      @     �W@      &@     �Z@      F@      @             �A@      B@              @     �E@      �?      2@      @     �I@      =@      @              &@      2@               @      ,@      �?      *@      @      8@      1@                      8@      2@               @      =@              @      @      ;@      (@      @              .@     �@@                      *@      @     @S@      @     �K@      .@      �?                       @                      @       @      4@      �?      "@       @      �?              .@      ?@                      @       @     �L@      @      G@      *@              4@     `k@     pw@      @@      J@     pt@     �T@      �@      e@     p@     �q@      9@      @     �O@     @d@      (@      (@     �]@      .@     �w@      N@     `m@     @Z@      @       @      &@     �H@      @       @      8@      �?     �c@      ,@      U@      8@               @      $@      @@      @       @      .@      �?      I@      *@      D@      0@                      �?      1@                      "@              [@      �?      F@       @              �?      J@     @\@       @      $@     �W@      ,@     �k@      G@     �b@     @T@      @      �?      D@     �S@      @      @     �T@      ,@     �\@      E@     �R@      O@      @              (@     �A@      @      @      *@              [@      @      S@      3@              1@     �c@     �j@      4@      D@      j@      Q@     0p@      [@     �p@     �f@      3@      .@     �\@      a@      .@     �A@     `a@      L@     �W@     @V@     �^@     �\@      0@      @     �P@     @S@      (@      ;@      Y@      6@      O@     �H@      U@      L@       @      &@      H@      N@      @       @     �C@      A@     �@@      D@      C@     �M@       @       @      E@      S@      @      @     @Q@      (@     �d@      3@     @b@     �P@      @       @      =@     �I@      @             �@@      $@     @\@      @     �X@      @@      @              *@      9@       @      @      B@       @     �I@      0@     �G@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ5�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @%��O}@�	           ��@       	                   �5@l��@	@�           ��@                           �?���C��@�           ��@                           �?|�&C�@S           ��@������������������������       ��K��:�@U            �a@������������������������       �a6� @�            Px@                           @���~��@�           X�@������������������������       �u��&�@�           ��@������������������������       ����g/@             :@
                           �?�o���@�           ��@                           �?}{:�@�            �s@������������������������       ���`x�@Y            �`@������������������������       �	����@v            �f@                           �?����k	@'           @�@������������������������       �;��
��
@�            �u@������������������������       ��.˛(�@F           ��@                           �?mH�Z�c@�           �@                           �?q�����	@�           �@                          �?@��yL�
@�            @q@������������������������       �ӛ��/�	@�             p@������������������������       �.Q���" @	             2@                           @$����@           �z@������������������������       �r$(֭�@�            @x@������������������������       ���_x��@            �B@                           �?�%c�J,@           �{@                           @�"m@�G @R             a@������������������������       ��3:�BP@#            �M@������������������������       �u���?/            @S@                           @\���3@�            ps@������������������������       �%ԩn[+@O            �_@������������������������       ����RzP@u             g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     @r@     0�@      8@     �O@      {@     �W@     0�@     �n@     x�@     pu@      >@      $@      i@      z@      "@     �C@     `r@     �O@     8�@     �e@     ��@     �l@      7@              S@      n@       @      2@      a@      *@     ��@     @S@     �v@     �\@      @              2@     �U@              @      9@       @     �m@      0@     �\@      <@      �?               @      <@               @      &@              @@      &@     �B@      &@      �?              $@      M@              �?      ,@       @     �i@      @     �S@      1@                      M@     `c@       @      .@     �[@      &@     �r@     �N@     �n@     �U@      @              L@     �b@       @      &@     �[@      "@     Pr@      N@     `n@     @T@      @               @      @              @               @      @      �?       @      @       @      $@     @_@     �e@      @      5@     �c@      I@     @j@      X@     �i@     �\@      1@              A@     �F@      �?      @      @@      @     @T@      ,@     �O@      C@      @              5@      4@              @      2@      �?      0@       @      :@      8@      @              *@      9@      �?              ,@       @     @P@      (@     �B@      ,@              $@     �V@     @`@      @      2@     �_@     �G@      `@     �T@     �a@      S@      ,@       @      ?@      J@      @      $@     �H@      <@      =@     �K@     �@@      @@      *@       @      N@     �S@       @       @     @S@      3@      Y@      ;@     �[@      F@      �?      .@     �V@     �d@      .@      8@     �a@      ?@     �o@      R@      k@     �\@      @      .@      R@     �Y@      ,@      1@      Y@      >@     �W@      L@     @\@     �S@      @       @      >@      B@      &@      $@      ?@      2@      C@      2@     �B@     �B@       @              :@      A@      &@      "@      <@      2@      C@      2@     �B@     �B@       @       @      @       @              �?      @                                                      @      E@     �P@      @      @     @Q@      (@     �L@      C@      S@      E@      @      @     �C@     �N@      @      @     �P@      "@     �G@     �@@     �R@      D@      @      @      @      @              �?       @      @      $@      @      �?       @                      3@     �O@      �?      @      D@      �?      d@      0@      Z@      B@                      @      "@              �?       @             �N@             �E@       @                      @      @                      @              <@              &@      @                      �?      @              �?      @             �@@              @@      @                      *@      K@      �?      @      @@      �?     �X@      0@     �N@      <@                      @      ?@              @       @             �B@      *@      0@      (@                      @      7@      �?      @      8@      �?      O@      @     �F@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�"�^/@�	           ��@       	                    �?�^�8X�@�           ��@                           �?�5�]�3	@S           P�@                           �?]�G�@�            �r@������������������������       �����@W            �b@������������������������       �B3-p<�@]            `b@                           @q�(��	@�           �@������������������������       �7�����	@�           8�@������������������������       �9K˕}�@             :@
                           @W����@t           �@                           �?���b��@	           �z@������������������������       ��P혀]@W            �`@������������������������       �DY� ��@�            pr@                          �4@�#A���@k           T�@������������������������       ��4����@�           (�@������������������������       �(:`NŮ@�           ��@                          �2@����v�@�           ��@                           �?��� @�             s@                          �0@$$g��?P             ^@������������������������       ��A�c�)�?             2@������������������������       �^��p��?D            �Y@                          �1@��􋹒@s             g@������������������������       �'ϲ��@<             W@������������������������       �`ţ8��@7             W@                           @�G�ٔ@           p�@                           �?+�R��R	@�           �@������������������������       �H�F%_�@q            @g@������������������������       ��ʷ�n�	@,           0|@                           @$15i��@}             j@������������������������       �M��@r            �g@������������������������       ��Ъ��@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      q@     �@      9@     �I@     �{@     �S@     ��@     �j@     ��@     0x@      B@      "@     @e@     �w@      .@      A@     `s@      L@     �@      b@     �@     �p@      =@      "@     @X@     �`@      (@      *@     �a@      ;@     @b@     �X@     �c@     �]@      3@              9@      H@      �?              D@       @      P@      1@     �Q@      ;@       @              (@      *@                      9@              D@      @      D@      1@                      *@     �A@      �?              .@       @      8@      ,@      ?@      $@       @      "@      R@      U@      &@      *@     @Y@      9@     �T@     �T@     @U@      W@      1@      @     �P@      U@      &@      *@     �X@      9@     �T@     �R@      U@      V@      *@       @      @                               @                      @      �?      @      @             @R@     `o@      @      5@      e@      =@     ��@      G@     |@     �b@      $@              7@     �L@              @     �K@      *@      Y@      6@      Y@      H@      @               @      &@              �?       @      @     �G@      �?      E@      &@      �?              .@      G@              @     �G@      $@     �J@      5@      M@     �B@       @              I@     @h@      @      ,@     �\@      0@     �~@      8@     �u@     �Y@      @              2@      W@      �?      "@     �@@      @     `u@      "@     @f@     �K@                      @@     �Y@       @      @     @T@      (@     �b@      .@     `e@     �G@      @      "@     �Y@     �d@      $@      1@      a@      6@     Pq@     @Q@     @k@     �]@      @      �?      3@      B@              �?      ;@             �[@      (@      Q@      =@                      @      @                      "@             @Q@       @      6@      $@                              �?                      @               @              @      �?                      @      @                      @             �N@       @      2@      "@              �?      .@      @@              �?      2@              E@      $@      G@      3@                      @      0@                      @              @@      @      3@      "@              �?      &@      0@              �?      *@              $@      @      ;@      $@               @     �T@      `@      $@      0@     �[@      6@     �d@     �L@     �b@     @V@      @       @     �R@     �Z@      $@      ,@     �V@      5@     �T@      J@     @Y@      R@      @              :@      >@              @      8@              B@      *@     �A@      3@               @      H@      S@      $@      &@     �P@      5@     �G@     �C@     �P@     �J@      @              "@      6@               @      4@      �?     �T@      @     �H@      1@      �?              @      2@               @      0@      �?      T@      @     �F@      1@                      @      @                      @              @              @              �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJz
 hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?U ��wQ@�	           ��@       	                   �;@d�M]	@�           ��@                           �?���p�	@W           �@                           �?������@           py@������������������������       ��N�
@k             e@������������������������       �� F'�@�            �m@                          �4@�{���	@S            �@������������������������       �!=u)y�@           @y@������������������������       �}�OM�	@O           ��@
                           �?P>�H)	@�            0p@                           @�׼�^Z@>            @\@������������������������       ����-�F@/            �U@������������������������       ���X�@             ;@                          �<@���g�@e            @b@������������������������       ��0+�4	@             ?@������������������������       ���Ȱ�@P            �\@                          �4@�!P���@�           �@                           �?���d�@�           �@                           @���Y�&�?           �|@������������������������       ����j�@:            �W@������������������������       ��PP��7�?�            �v@                           �?/�R+@�           ��@������������������������       �p~$0��@            �J@������������������������       �$�L�@�           �@                           @����@�            �@                           �?��ɒ�L@�           ��@������������������������       �6�\t�@?           @@������������������������       �R� �@H           h�@                            �?Q���y�@            �C@������������������������       ��|J��@
             4@������������������������       �\���Q.�?             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     h�@      ?@     �J@     �z@      W@     ��@     �l@     ȉ@     �v@      ?@      .@     �c@     `m@      5@      =@      n@     �N@     �l@     �b@     �o@     �f@      9@      $@     @_@     @h@      *@      8@      i@     �G@      k@      _@     �l@     �`@      9@              C@     @Q@      @      @      G@      @     �X@      5@      V@      =@      @              ,@      =@                      .@              H@      @      G@      &@      �?              8@      D@      @      @      ?@      @     �I@      1@      E@      2@      @      $@     �U@     @_@      $@      4@     @c@     �D@     @]@     �Y@     �a@     �Y@      5@      @      C@      B@      @      @     @R@      ,@     �P@     �B@     �P@      J@       @      @     �H@     @V@      @      0@     @T@      ;@      I@     �P@     �R@     �I@      *@      @      @@     �D@       @      @      D@      ,@      ,@      8@      9@     �I@              �?       @      :@      @      @      1@      &@      @      $@      $@      5@                      @      :@      @      @       @      $@      @      @      @      1@              �?      @                              "@      �?              @      @      @              @      8@      .@      @       @      7@      @      &@      ,@      .@      >@              @      @       @      @      �?      @      �?      @               @      @                      3@      *@       @      �?      2@       @       @      ,@      *@      9@              @     �a@      r@      $@      8@     @g@      ?@     Ȉ@     �T@     ؁@      f@      @              H@     �c@      @      (@     �Q@      @     �@      =@     �r@     �U@                      1@     �D@               @      3@              o@      @     @Z@      6@                      @      @                       @              B@              <@      $@                      &@      A@               @      &@             �j@      @     @S@      (@                      ?@     @]@      @      $@     �I@      @     Pp@      9@      h@      P@                              "@              @       @      @      (@      @       @      @                      ?@      [@      @      @     �E@              o@      4@      g@     �N@              @     @W@     �`@      @      (@      ]@      <@     �q@      K@     q@     �V@      @      @     @T@     �`@      �?      (@     �[@      9@     �q@      G@     �p@     �V@      @      @      <@     �N@              @     �N@      $@     �a@      .@     �`@     �B@      @             �J@     �Q@      �?      @     �H@      .@     �a@      ?@     �`@      K@      @              (@              @              @      @      @       @      @                              @              @              �?      @      �?      @      @                              @                              @               @      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�x�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @w�l�3@�	           ��@       	                    �?�>�5��@d           &�@                          �;@;����@�           �@                           �?;�4�՛@M           P�@������������������������       �,����@           `y@������������������������       ��d��	@I           ��@                           @k�4��@�             n@������������������������       ��z��2A@s            �e@������������������������       ���e�L@+            �P@
                           �?@=�7�@y           p�@                            �?@f{�@o            `e@������������������������       ���@��@'             M@������������������������       ���I�@H            @\@                          �4@	�3F<[@
           0z@������������������������       �u/ �H�@w            �f@������������������������       �K����@�            �m@                          �7@��I7@F           ؚ@                           �?3��u�;@O           ��@                           @X�KS@3           P}@������������������������       �4����?�            �t@������������������������       ��.�;�@a             a@                           @���A)@           ؊@������������������������       ��5���@�           �@������������������������       ��Ғ�Z�@�            @k@                           @"��� .@�            `x@                           @�bluf?@�            �k@������������������������       �;��uA�@=            �W@������������������������       �ʅT�`�@T            �_@                            �??��4Z%@f             e@������������������������       �!���oB@             D@������������������������       �'`�!H@N             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     pr@     X�@      >@      H@     �}@     �R@      �@     `j@     @�@     �w@     �A@      &@     `j@      s@      3@      B@     �u@     �J@     �v@     �e@     �x@     �o@      <@      &@     `c@     �j@      2@      >@     0q@      C@     @k@     �`@     pq@     �i@      <@       @      `@     �g@      (@      9@     �m@      :@     �i@     �[@      p@     �a@      9@             �C@      L@      @      @      L@      �?     �T@      8@     @Z@      >@      @       @     �V@     �`@      @      5@     �f@      9@      _@     �U@     �b@      \@      5@      @      :@      ;@      @      @      C@      (@      (@      6@      7@      P@      @      �?      5@      8@      @      @      5@       @      @      .@      0@     �I@       @       @      @      @              �?      1@      @      @      @      @      *@      �?              L@     �V@      �?      @     �Q@      .@      b@     �D@     �]@     �G@                      .@      (@              �?      0@       @      N@      @     �H@      "@                      @      @              �?      @      �?      3@              7@       @                      (@      @                      (@      �?     �D@      @      :@      @                     �D@     �S@      �?      @      K@      *@      U@      A@     �Q@      C@                      @     �B@      �?      �?      7@      �?      N@      $@      ?@      ,@                     �B@      E@              @      ?@      (@      8@      8@     �C@      8@              �?      U@      o@      &@      (@     �_@      5@     Ѓ@      C@     �y@      _@      @             �N@     `j@      $@       @     �R@      0@     �@      4@     0s@     �R@      @              ,@     @R@      �?       @      5@      @     �m@       @     �V@      .@       @              @     �H@                      *@      @     �f@      @     �P@      "@                      "@      8@      �?       @       @              L@      @      9@      @       @             �G@     @a@      "@      @      K@      (@     �r@      (@      k@     �M@      @              ?@      Y@      @      @     �A@      @     @o@      @      e@     �@@      @              0@      C@      @       @      3@      @     �J@      @     �G@      :@              �?      7@      C@      �?      @      J@      @     @W@      2@     �Y@      I@       @      �?      0@      ;@              @      =@      �?     �L@      @     @P@      .@       @      �?      $@      @              �?      .@              :@      �?      ?@      @                      @      5@               @      ,@      �?      ?@      @      A@      &@       @              @      &@      �?      �?      7@      @      B@      *@      C@     �A@                       @       @                      @      @      &@      @      @      @                      @      "@      �?      �?      4@              9@       @      @@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ�5HhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�e�x1@�	           ��@       	                     �?I���@�           X�@                           �?j�G�@�            �v@                           @�)��V@c             c@������������������������       ��if;@2            �S@������������������������       �eŅ-��?1            �R@                           �?[?�@}            �j@������������������������       �ة�t#@.            �U@������������������������       ��������?O            �_@
                           @Ԍ�H
@�           ��@                           �?���1�@O           `�@������������������������       ��9�L>�@�             j@������������������������       ���(�@�            �u@                           @�N���@h           �@������������������������       �m��*X @�            �r@������������������������       �DS��g@�            Pq@                           �?#��O.@           �@                           �?�4@�@�           ȅ@                          �;@rC�Ӑ@�             t@������������������������       ����9�@�             p@������������������������       �(�߾�@%             P@                           @|U2&6@�            �w@������������������������       ��y��Ĥ@f            �b@������������������������       ����.ܛ@�            @l@                            �?������@h           �@                           @|}i*	@;           �~@������������������������       ��6�	@L            �_@������������������������       ��1��s@�             w@                           @��祔@-           0�@������������������������       ��p,uh	@�           ��@������������������������       �M�()��@G           �~@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �s@     ��@      5@     �N@     P|@     �R@     �@      h@     �@      x@     �@@      @     �S@     �g@      @      (@     @a@      $@     `�@     @P@     0u@     �^@      @              &@      I@              �?      8@      @     �b@      7@      T@      2@      @              �?      *@              �?      0@      @     �P@      "@     �@@      @      @              �?      "@                      (@      @      4@      "@      1@      @      @                      @              �?      @              G@              0@      @                      $@     �B@                       @             �T@      ,@     �G@      (@       @              @      $@                      @              0@      *@      7@       @       @              @      ;@                      �?             �P@      �?      8@      @              @      Q@     �a@      @      &@     �\@      @     pw@      E@     0p@      Z@              @     �B@      U@      @      "@     �S@      @      a@      ?@      W@     �R@                      (@      A@                      9@       @      P@      @      D@      9@              @      9@      I@      @      "@      K@      @      R@      9@      J@     �H@                      ?@     �L@               @     �A@      �?     �m@      &@     �d@      >@                      0@      8@              �?      2@             �c@      "@     @P@      @                      .@     �@@              �?      1@      �?     �T@       @     �Y@      7@              $@     �m@     �w@      0@     �H@     �s@      P@     P}@     �_@     �|@     `p@      ;@             �O@      \@       @      $@     �Q@      @     �g@      8@     �c@     �L@      @              I@     �L@       @       @      @@      @     �I@      (@     �N@      D@      @              E@      F@       @      @      :@              G@      &@      L@      6@      @               @      *@              @      @      @      @      �?      @      2@                      *@     �K@               @     �C@      @     `a@      (@     @X@      1@                      &@      0@               @      6@       @     �J@      @      @@       @                       @     �C@                      1@      �?     �U@      @     @P@      "@              $@     �e@     �p@      ,@     �C@     �n@      M@     pq@     �Y@      s@     �i@      7@      �?     �P@      T@      @      ,@      O@      (@     �S@      B@     @Q@      N@      $@              &@      0@              @      7@      @       @      ,@      4@      2@      @      �?      L@      P@      @      "@     �C@      @     �Q@      6@     �H@      E@      @      "@     �Z@     �g@      "@      9@     �f@      G@      i@     �P@     `m@      b@      *@      @      T@     �]@      @      ,@     @]@      A@      S@     �J@      _@      X@      &@       @      ;@     �Q@      @      &@     @P@      (@     @_@      ,@     �[@     �H@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�)%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�[BvN@�	           ��@       	                    @O�e�e@S           �@                           �?YPd�@�           ��@                          �2@�v`U@�            �v@������������������������       �u{�k�@o            `e@������������������������       ��`k��8@�            `h@                           �?���iE\@�           �@������������������������       �'J?ٹ@/           `@������������������������       �CQFC/@x            �h@
                           �?���~@D@�           ��@                          �3@��"f��?           `z@������������������������       �%��F�?�            @s@������������������������       ���Bq�?@            �\@                           �?�4Ʉ�@�           ��@������������������������       ����@             G@������������������������       ���V��@�           p�@                          �<@��!P2�@;           �@                           @��)�:}@d           p�@                          �;@����H�@U           Ќ@������������������������       ��}7�ω@%           ��@������������������������       �]7�@0             Q@                           �?	�~��T	@            |@������������������������       �q�aa�	@s            @g@������������������������       ��=��@�            �p@                           @nu'Q�}	@�             v@                            �?�6��L�	@X            @b@������������������������       �G�[g��@+            �P@������������������������       ��-�'	@-            �S@                           @!��<�P@            �i@������������������������       ����r��@`            �b@������������������������       � ;O���@            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     �p@     ��@     �B@      D@     p@      S@      �@     �i@     �@     pv@      B@      @     �W@      t@      2@      2@     �m@      :@     ��@     �T@     8�@     �c@      (@      @      O@     �c@      &@      *@     �c@      2@     �l@      R@      l@     @[@      @       @      2@      O@      @      @     �P@       @      U@      <@      N@      :@      �?              @      @@      �?              E@       @      I@      "@      .@      ,@      �?       @      *@      >@      @      @      9@      @      A@      3@     �F@      (@              @      F@      X@      @      $@     �V@      $@      b@      F@     �d@     �T@      @      @      C@     @P@      �?       @     �R@      "@     �S@      @@     �^@     �O@      @              @      ?@      @       @      1@      �?     @P@      (@      E@      4@                      @@     �d@      @      @     �S@       @     @}@      &@     `r@      I@      @              (@     @P@                      .@             �k@      @      X@      "@      �?              $@      B@                      &@              d@      @     @S@      "@      �?               @      =@                      @              N@              3@                              4@     �X@      @      @     �O@       @      o@      @     �h@     �D@      @              �?      "@                      (@      @      @       @      &@                              3@     �V@      @      @     �I@       @     `n@      @     `g@     �D@      @      6@     �e@      n@      3@      6@     �p@      I@     �r@      _@     �q@      i@      8@      0@      a@     �g@      (@      .@      l@     �B@     �p@     @V@     �m@      `@      4@      "@     �U@     ``@      @      @     `b@      >@     �i@      D@      e@     �T@      &@      @      U@      ]@      @      @     �a@      =@     �g@      B@     �c@      S@      $@      @      @      .@              �?      @      �?      ,@      @      (@      @      �?      @     �H@     �M@      @      $@     @S@      @     �N@     �H@     �Q@      G@      "@      @      (@      =@      @      @      B@      @      ,@     �@@      1@      4@      @             �B@      >@      @      @     �D@      @     �G@      0@     �J@      :@      @      @     �B@      I@      @      @     �E@      *@      A@     �A@      F@      R@      @      @      "@      5@      @      @      ,@      @      (@      1@      5@      >@       @               @      @              @      @      @      @      $@       @      5@       @      @      @      .@      @      �?      "@              @      @      *@      "@                      <@      =@      �?       @      =@      $@      6@      2@      7@      E@       @              1@      :@      �?       @      1@      $@      (@      2@      .@      ?@       @              &@      @                      (@              $@               @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ`K�9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?@�1�5@�	           ��@       	                   �8@v�r �@           �@                           �?�ds�@z           �@                           �?V@����@B           `@������������������������       �~�ͯ��@_            �a@������������������������       �Q�3U)?�?�            pv@                            @ÿ�1@8           �~@������������������������       �Cr��i@�            @v@������������������������       ��/|%�L@U            �`@
                           �?H|���@�            �l@                            �?XÇ,�g@Z             a@������������������������       �2�^m?r@3            �R@������������������������       �_(ٜU@'             O@                          �>@�`X�@F@A            @W@������������������������       �9��~2d@9             U@������������������������       �//�jsx @             "@                          �4@�y��@�           �@                          �1@��J[~�@�           ��@                           �?��Z1��@�            �v@������������������������       �8P3[9�@>             [@������������������������       �B^1��R@�            �o@                            �?O��C�@�           �@������������������������       ���rkTX@             h@������������������������       �E���#@~           �@                           �?}nm���@�           \�@                           �?��q�s@J             ]@������������������������       ��H>W��@             A@������������������������       ��l��@3            �T@                           @���@x           ��@������������������������       �u�E@|           ��@������������������������       �D�已x@�           `�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �p@     ��@     �@@     �H@     P}@     �R@     ��@      l@      �@     pu@      ?@      @      S@     �b@      @      @      Y@      @     �~@      E@     �p@     @R@       @              M@     �]@      @       @      R@      �?     �{@      :@     @k@     �E@      @              6@     �N@      �?      �?      C@      �?     �o@      *@     @V@      3@      @              @      6@      �?              1@             �G@      @      >@      $@      @              0@     �C@              �?      5@      �?     �i@      @     �M@      "@                      B@     �L@       @      �?      A@             �g@      *@      `@      8@      @              9@     �E@       @              9@             �b@      @     �V@      (@      @              &@      ,@              �?      "@              E@       @      C@      (@              @      2@      ?@              @      <@      @      G@      0@      G@      >@      �?      @      2@      6@              @      4@      �?      *@      &@      4@      7@      �?      @      @      .@              �?      @      �?      @      @      &@      4@      �?              (@      @               @      .@              @       @      "@      @                              "@                       @      @     �@@      @      :@      @                              "@                      @      @      @@      @      9@      @                                                      @              �?      �?      �?       @              ,@      h@     �y@      >@      F@     w@      Q@     �@     �f@     �@     �p@      7@      @     �K@      c@      &@      0@     �`@      3@     �u@     @S@     �o@     �\@      &@              $@     �F@              @      B@      @     �`@      0@     @U@      <@                       @      &@              �?      0@      @      2@       @      <@      .@                       @      A@               @      4@             @]@       @     �L@      *@              @     �F@      [@      &@      *@     �X@      0@     �j@     �N@     �d@     �U@      &@              $@      2@                      6@      @     @Q@      1@     �A@      0@      @      @     �A@     �V@      &@      *@      S@      *@     @b@      F@     �`@     �Q@       @      &@      a@     0p@      3@      <@     `m@     �H@     �l@     �Z@      p@     `c@      (@      @      *@      2@              "@      8@      @      @      $@      8@      @      �?      �?       @      $@                      @      �?                       @       @      �?       @      @       @              "@      5@      @      @      $@      0@      @               @      _@      n@      3@      3@     `j@     �F@     �k@      X@      m@     �b@      &@      @     �F@     �Y@      *@      @     �V@      :@     @\@     �@@     �U@      T@              @     �S@     `a@      @      *@     @^@      3@     �[@     �O@      b@     �Q@      &@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJoV�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���υN@�	           ��@       	                    �?���ƪ�@v           `�@                           �?��8�l�@�           ��@                          �;@�w�.[@�            pr@������������������������       �iX����@�            �p@������������������������       �e���ƶ@             >@                           �?��߾\@�            �u@������������������������       ��h��2�@�            �n@������������������������       ��|e�@:            �X@
                          �6@G���(`	@�           Ę@                           �?-�i@/           �@������������������������       �jZ���@�           Ѓ@������������������������       �9|���@�            �p@                           �?)U�	
@�           p�@������������������������       �ȃ&��@k            �d@������������������������       �N��h*
@A           H�@                            @�U��@            d�@                           �?���s9@u           �@                            �? 
τ�T@'           ~@������������������������       �x��T���?P            �]@������������������������       �x0�嫯@�            �v@                          �6@��n�,�@N            �@������������������������       �WV�m$@�           ��@������������������������       �����@�            �r@                           @ĥ��F�@�            �q@                           @W75L�E�?\            @c@������������������������       ��]ղ���?*            �S@������������������������       ��8<XJ��?2             S@                           �?qW�d*@O            �_@������������������������       �$nX�/�@)            @Q@������������������������       �[6<�R�@&            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      s@     `�@      ;@     �I@     �{@     @S@     P�@     @o@     ؈@     0t@      B@      0@     @l@     @u@      2@      B@     @s@      M@     �w@     �i@     �w@      l@      @@       @     �P@     @U@      �?      @      Q@      @     �f@      <@      b@      J@       @       @      :@     �D@      �?      @      C@      @     �V@      &@     �K@      7@                      7@     �A@      �?       @      B@       @     �V@       @     �I@      1@               @      @      @               @       @      �?      �?      @      @      @                     �D@      F@              �?      >@      �?     @V@      1@     �V@      =@       @              @@      C@              �?      9@             �L@      1@      J@      8@                      "@      @                      @      �?      @@              C@      @       @      ,@     �c@     �o@      1@      ?@      n@      K@      i@      f@     �m@     �e@      >@      $@     �R@     `d@      @      ,@     �b@      4@     �a@     @V@     �`@     �V@       @      $@     �N@     �[@      @      $@     @[@      0@     �T@      N@      X@      Q@       @              *@     �J@      �?      @      E@      @     �M@      =@      C@      6@              @     @U@      W@      *@      1@     @V@      A@      M@     �U@     �Y@     �T@      6@      �?      $@      =@      �?       @      2@      @      3@      5@      @@      3@      @      @     �R@     �O@      (@      .@     �Q@      <@     �C@     �P@     �Q@      P@      .@      �?      T@      o@      "@      .@     �`@      3@     p�@      G@     �y@     �X@      @      �?     �Q@     @l@      @      "@     @\@      2@     �@      D@     @t@     @U@      @              .@     @T@       @             �@@      "@     @k@      "@     @V@      9@                              &@       @              &@       @     @Q@       @      1@      @                      .@     �Q@                      6@      @     �b@      @      R@      4@              �?      L@      b@      @      "@      T@      "@     pr@      ?@     `m@      N@      @              =@     �X@      @      �?      E@      @     �m@      @      d@      C@      @      �?      ;@      G@      �?       @      C@      @      M@      8@     �R@      6@                      "@      6@      @      @      4@      �?     @[@      @     �V@      *@      �?              @      *@                      "@      �?     @Q@             �K@      �?      �?               @      "@                              �?     �C@              ;@                              @      @                      "@              >@              <@      �?      �?              @      "@      @      @      &@              D@      @     �A@      (@                              @      �?      @      �?              7@       @      :@       @                      @      @       @       @      $@              1@      @      "@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�8���[@�	           ��@       	                    �?2��	��@z           n�@                           �?��C+,	@           �@                           @�+���	@z           Ȃ@������������������������       ��%ޚJ�@�            �v@������������������������       �HgG�8�@�            �m@                           �?L}Rw�@�           ��@������������������������       �m�6�|�@�            pw@������������������������       ���&�3	@�           X�@
                           �?���|MF@w           ��@                          �9@�@<x@n            `e@������������������������       ������@]            `b@������������������������       �.�X��k@             8@                          �5@�3m��/@	           y@������������������������       �6��	U�@�            @k@������������������������       ����*j@}            �f@                            �?l>8 �@/           H�@                          �7@��[c@[           p�@                           @�H>0�@�           (�@������������������������       �����@X           ��@������������������������       ��B燁5@�            �i@                           �?}�j�ϳ@�             i@������������������������       �*r�1V�@>            @Y@������������������������       �t�D�r�@D             Y@                          �4@�H!X�@�            �@                           �?7���2@�            `w@������������������������       ����]:��?f             c@������������������������       �Y��{�@�            �k@                           @���»d@�            �v@������������������������       �!{Ǩ�Z@�             t@������������������������       ���4��@             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     0�@      =@     �M@      |@      U@      �@      k@     H�@     �w@      @@      *@     �m@      t@      4@     �I@     �s@      P@     �v@     �e@     �w@     �p@      8@      *@     �g@     `o@      2@      E@     @o@     �H@     �l@     �_@     0p@     @j@      6@       @     �P@     @[@      &@      8@      V@      2@     �S@     �L@      M@      T@      $@       @     �C@     @P@      $@      *@     �L@      0@      O@      2@      B@     �G@                      ;@      F@      �?      &@      ?@       @      0@     �C@      6@     �@@      $@      &@     �^@     �a@      @      2@     @d@      ?@      c@     @Q@      i@     @`@      (@              ?@      N@       @      @      H@      �?     @Q@      6@     �R@     �M@       @      &@     �V@     �T@      @      (@     �\@      >@      U@     �G@     �_@     �Q@      $@              H@     �Q@       @      "@      Q@      .@     �`@      G@      _@      K@       @              0@      &@                      ,@      �?     @Q@      @      H@       @      �?              .@      @                      &@      �?     �P@       @      B@       @                      �?      @                      @               @      �?      (@              �?              @@      N@       @      "@      K@      ,@      P@     �E@      S@      G@      �?              @      >@       @      @      9@      @      H@      4@     �H@      <@                      9@      >@              @      =@      $@      0@      7@      ;@      2@      �?      @     @T@     �h@      "@       @     �`@      4@     ��@     �F@     �x@     �]@       @             �E@      _@      @      @      P@      0@     pv@      9@      l@     �R@      �?              7@     @Z@      @      @      I@      &@     ps@      &@     @e@      H@      �?              ,@      R@      @              =@      @     @o@      @     �\@     �C@      �?              "@     �@@       @      @      5@      @     �N@      @      L@      "@                      4@      3@                      ,@      @      H@      ,@      K@      ;@                      .@      &@                       @              :@      @      9@      *@                      @       @                      @      @      6@      &@      =@      ,@              @      C@      R@      @       @      Q@      @     Ps@      4@     @e@     �E@      @              3@     �A@      @              2@              g@      $@     @V@      .@      �?               @      *@                      @              W@       @     �B@       @      �?              1@      6@      @              ,@              W@       @      J@      *@              @      3@     �B@      �?       @      I@      @     @_@      $@     @T@      <@      @      @      (@      @@      �?       @      B@      @     @]@       @     @S@      <@                      @      @                      ,@               @       @      @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ �rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?_=�AJ@�	           ��@       	                    @� 2@�           Ȑ@                           �?�Ƿ�-�@�           ��@                          �:@0#��G�@�            p@������������������������       ���s��(@�            �j@������������������������       �1~�5O�@             F@                           �?_S�1Pk@           `y@������������������������       �5�CP�@F            �Z@������������������������       �R�X	@�            �r@
                           @���pip@�            �y@                           �?*ʨ��|@�            0w@������������������������       �"׻;�F�?V            �_@������������������������       �B}
k�,@�            �n@                          �3@��)�@             D@������������������������       ���\�O� @	             .@������������������������       ���J��D@             9@                           �?���E@           .�@                            �?�i���@B           X�@                          �<@[��X�g@�            �t@������������������������       �6�+�ύ@�            �r@������������������������       �p�U~9 @             >@                            @WE{W��@g           ��@������������������������       �l�Z>5�@�            `k@������������������������       ���8_]�@�            @v@                           �?�`��}@�           0�@                          �1@<�ǔQ@�           ��@������������������������       ��Mݰ��@E            @Z@������������������������       �a}"g�@�           P�@                          �:@��ƻ �@�           d�@������������������������       �~�7�%@u           ��@������������������������       ��ʡ��@}             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     �@      8@      F@     �z@     �W@     ȏ@      m@     8�@     `w@      ?@      @     �R@     �a@      @      &@      _@      >@     ps@      U@     �g@     �U@      $@      @     �M@     �X@      @      "@     �Y@      :@      ]@     @R@     @[@      K@      $@       @      4@     �D@      �?      @      G@      "@     �D@     �B@      @@      2@      @              3@      B@      �?      @     �B@      @      D@      =@      7@      .@      @       @      �?      @                      "@      @      �?       @      "@      @               @     �C@     �L@       @      @      L@      1@     �R@      B@     @S@      B@      @               @      :@                      "@              6@      @      B@       @      �?       @      ?@      ?@       @      @     �G@      1@     �J@     �@@     �D@      A@      @              .@     �F@      @       @      6@      @     `h@      &@     �T@      @@                      ,@      E@                      6@      @     �f@      @     @S@      8@                              ,@                      @      @     �Q@              9@      "@                      ,@      <@                      0@      �?     �[@      @      J@      .@                      �?      @      @       @                      ,@      @      @       @                               @               @                      @              �?      @                      �?      �?      @                               @      @      @      @              ,@     @l@     @{@      2@     �@@     �r@      P@     �@     �b@     @�@      r@      5@              Q@      a@      @       @      O@      @      u@      C@      g@     �O@       @              ?@      L@      �?      @      2@      �?     �Y@      ,@     @Q@      A@       @              =@      K@      �?       @      2@      �?     �X@      "@     @Q@      2@       @               @       @               @                      @      @              0@                     �B@      T@       @      @      F@      @     @m@      8@      ]@      =@                      $@      <@                      2@      @     �U@      @     �L@      $@                      ;@      J@       @      @      :@             �b@      3@     �M@      3@              ,@     �c@     �r@      .@      9@     �m@      M@      w@     �[@     �x@      l@      3@      @      J@     �Y@      @      ,@      Z@      :@     �b@      @@      d@     @U@      *@              @      3@                      @              F@      @      4@      @              @      G@      U@      @      ,@     @X@      :@     �Z@      <@     �a@      T@      *@      @     �Z@     �h@       @      &@     �`@      @@     `k@     �S@     �m@     �a@      @      @     �P@      f@      @      @     �Z@      9@     �h@     @P@     `k@     �Y@      @      @     �C@      5@      @      @      =@      @      6@      *@      3@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���9�g@�	           ��@       	                    �?(^R��@s           N�@                           �?s)FGdQ	@�           X�@                          �;@��� �@+           @@������������������������       ��(�-3@           {@������������������������       �n�JO��@)            �P@                            �?E��7�	@�           ��@������������������������       �D�k*x	@�             u@������������������������       ���_6��	@�           ��@
                           �?|�1�E@}           ��@                            �?G^��'�@�             n@������������������������       �y�n*@+            �Q@������������������������       �<t4"=@n            @e@                            �?L�N��f@�            v@������������������������       ��?5�L@~            @h@������������������������       ��/��|@f            �c@                           @I@'�)@#           ��@                            @�	Ê*@�           T�@                          �4@�1 d�|@|           0�@������������������������       ���)@c           �@������������������������       ��n�͌@           �|@                          �3@�c�~10 @f            �e@������������������������       ��sU��6�?4            �V@������������������������       ��=�� @2             U@                          �7@Կ�r'�@A           h�@                           �?�߄�@�            pv@������������������������       ����s��@n            �e@������������������������       ���Tj-�@m             g@                           @v	�M�*@f            �d@������������������������       �6�V�@@            �Z@������������������������       ������@&            �M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �o@     p�@     �B@     �P@     �|@     �R@     ��@     @k@     ��@     Px@      >@      7@      f@     Pu@      =@     �H@     `s@     �L@     �w@     �f@      w@      q@      7@      7@     �b@     �n@      8@     �B@     �k@     �D@     �n@     �a@      p@     @k@      5@       @     �C@     �V@      @      @      O@      �?     �\@      =@     �X@      J@       @              @@     @S@      @      @      I@      �?     �Z@      :@     @X@      @@       @       @      @      *@              �?      (@              @      @       @      4@              5@     �[@     `c@      5@      >@     �c@      D@     �`@     �[@     �c@     �d@      3@       @     �A@      E@      �?      "@     �E@      1@     �J@     �E@      H@      B@      @      3@     �R@     @\@      4@      5@     �\@      7@     �S@      Q@     �[@     @`@      (@              ;@      X@      @      (@     �V@      0@      a@      E@      \@      K@       @              "@      <@      �?      @      G@       @     �M@      *@     �H@      5@      �?                      "@                      1@       @      1@       @      1@      @      �?              "@      3@      �?      @      =@      @      E@      &@      @@      0@                      2@      Q@      @      @      F@       @     �S@      =@     �O@     �@@      �?               @      ?@      @      @      .@      @     �H@      ,@      F@      1@      �?              $@     �B@              �?      =@      @      =@      .@      3@      0@               @     �S@      k@       @      1@     �b@      2@     ��@      B@     z@     @]@      @       @     �I@     `c@              @      Y@      @     @}@      3@     �q@      T@      @       @      G@      b@              @     �T@      @     �x@      2@     �k@     �R@      @              7@     �Q@              �?      8@      �?     `p@      @     �]@     �@@               @      7@     �R@              @     �M@      @     @`@      &@     �Y@      E@      @              @      $@                      1@              S@      �?     �M@      @       @              @      $@                      �?              E@      �?      A@                               @                              0@              A@              9@      @       @              ;@      O@       @      (@     �H@      &@     �d@      1@      a@     �B@       @              1@     �E@       @      $@      <@      @     �`@      @     @U@      6@       @               @      4@      @       @      6@       @     �M@      @     �B@      (@                      "@      7@      @       @      @      @     �R@       @      H@      $@       @              $@      3@               @      5@      @      ?@      (@     �I@      .@                      @      1@               @      @       @      <@      @      @@      "@                      @       @                      0@      @      @      @      3@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�\�VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?	d�jC@�	           ��@       	                   �2@#[z5*	@           ș@                            @l6��0�@�            �s@                            �?"�.�N@r            �e@������������������������       �"5n��@>            �X@������������������������       ����U�@4            �R@                          �1@9uN4,@Z            �a@������������������������       ���g��_@/             R@������������������������       �3ظ��o@+            @Q@
                           �?|���	@F           ܔ@                           �?؝�pr
@�            �x@������������������������       �}a��B@q            �e@������������������������       �؁�*�@�             l@                           @(��
@S           H�@������������������������       ��FAJw"
@�             i@������������������������       ��X���	@�           �@                           �?�>�s��@�           ��@                           �?�B���@�           H�@                          �3@�a�� @            {@������������������������       ���*;�G�?}            �h@������������������������       �NBq�<�@�             m@                           @C����$@�            �u@������������������������       �O��2�� @�            �o@������������������������       �3�f@>            @W@                            �? d#���@�           8�@                          �2@���$��@           ��@������������������������       �"���Է@�             o@������������������������       �{i����@�            �@                          �4@)��F�@�           ��@������������������������       �����@�            pq@������������������������       ����_�@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �p@     ؁@      =@     �M@      }@      T@     8�@      i@     ��@     Pw@      ?@      3@     `b@     �o@      4@     �A@      p@     �I@      i@      _@      r@     �l@      9@              1@     �A@      �?      @      M@      @     �M@      5@     �S@      B@      @              @      9@                      A@      �?      ?@      .@      B@      6@      @              @      0@                      3@      �?      ,@      $@      ;@      @       @              @      "@                      .@              1@      @      "@      0@      �?              $@      $@      �?      @      8@      @      <@      @      E@      ,@                      @      @      �?      �?      &@              5@      @      0@      $@                      @      @               @      *@      @      @      @      :@      @              3@     @`@     `k@      3@      @@     �h@     �G@     �a@     �Y@     @j@     @h@      6@              F@     @Q@      �?      @     �O@      @     �H@      9@     �V@     �F@       @              4@      9@      �?      @      >@      @      2@      ,@      E@      2@                      8@      F@              @     �@@              ?@      &@     �H@      ;@       @      3@     �U@     �b@      2@      :@     �`@      F@     @W@     �S@     �]@     �b@      4@      $@      3@      6@      @      �?      ?@      *@      &@      3@     �D@      5@      @      "@     �P@      `@      (@      9@      Z@      ?@     �T@     �M@     �S@      `@      ,@      �?     �^@     �s@      "@      8@      j@      =@     ��@      S@     ��@     �a@      @              B@     @V@      �?      �?     �F@      @     Pv@      (@     @h@     �@@       @              7@      H@              �?      <@      �?      k@      @     �V@      4@                      *@      1@              �?       @              Z@       @      I@      @                      $@      ?@                      4@      �?      \@      @      D@      0@                      *@     �D@      �?              1@      @     �a@      @      Z@      *@       @              &@     �A@                      @      @     @[@      �?     �R@      @      �?               @      @      �?              $@              @@      @      =@      @      �?      �?     �U@     �l@       @      7@     `d@      6@     �y@      P@     �v@     �[@      @              L@     �]@      @      .@      T@      1@      m@      A@     �l@      Q@      �?              @     �A@      @       @      "@      �?     �Z@       @     �P@      2@                      J@     �T@      �?      *@     �Q@      0@     �_@      @@     `d@      I@      �?      �?      ?@     �[@      @       @     �T@      @      f@      >@     @a@      E@      @              $@      G@      �?      @      ;@       @      [@      "@      L@      .@              �?      5@      P@       @      @      L@      @      Q@      5@     �T@      ;@      @�t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?"���?@�	           ��@       	                   �3@6�I|�@7           �@                           �?�a�D��@�           ��@                            @��&���@x            @f@������������������������       �� ���@>            �X@������������������������       �������@:            �S@                          �1@�2��@2           �~@������������������������       ��8d�� @�            `l@������������������������       �e� ���@�            �p@
                          �8@e_P:�g@�           @�@                           @�F>z8�@�           H�@������������������������       �Ǭh��@�            0s@������������������������       ��r�'r@�            `u@                          �9@�Χ)�@�            �u@������������������������       ��˟��@*             R@������������������������       �M�W�Ų@�            pq@                          �7@�6�[@�           ��@                           �?�<)u[@�           p�@                            �?o��,��@           �|@������������������������       ��+��@�            �o@������������������������       �z����@�             j@                           �?ww-d�T@�           4�@������������������������       ��@r�8�@3            �U@������������������������       �����f@�           ��@                          �<@gY�[z�@�           0�@                           �?�L@/           �}@������������������������       ����@@             Z@������������������������       ���l4�@�            @w@                            �?Άo�M	@�            @i@������������������������       �l)]�Z@P            �\@������������������������       ��S��F@7            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     X�@      A@      K@     P~@     �S@     ��@     �g@     ��@     �v@      @@      @      `@      n@      5@      7@     �k@      B@     �}@     @P@     pr@     �b@      $@      �?      D@     @V@               @     �Q@      @     `p@      .@     �`@      I@       @      �?      (@      9@                      ?@      @      D@      @      =@      :@       @      �?      @      4@                      2@      @      .@      @      1@      &@       @              @      @                      *@       @      9@      �?      (@      .@                      <@      P@               @      D@             �k@       @     @Z@      8@                      @     �A@               @      2@             @^@      �?      B@      $@                      8@      =@                      6@             @Y@      @     @Q@      ,@              @      V@      c@      5@      5@      c@      ?@     �j@      I@      d@     �X@       @             �P@      W@      .@      ,@     �W@      2@     �d@      0@     �[@     �H@      @             �C@      K@      (@      &@      L@      @      G@      .@      B@      ;@      @              <@      C@      @      @     �C@      &@      ^@      �?     �R@      6@      @      @      5@      N@      @      @     �L@      *@     �H@      A@     �I@     �H@      �?              @      @      �?      �?      4@       @      @      (@       @      (@              @      ,@     �K@      @      @     �B@      &@     �F@      6@     �E@     �B@      �?      $@      g@     �s@      *@      ?@     `p@      E@     ��@     @_@     �~@     �j@      6@      @     �`@     @m@      @      0@     �b@      9@     �z@     �Q@     �v@     �^@      &@             �D@     �L@       @      �?      A@             `e@      @      `@      6@      �?              6@      >@       @              ,@             �W@             �S@      ,@                      3@      ;@              �?      4@              S@      @      I@       @      �?      @     �V@      f@      @      .@     �\@      9@      p@      P@     �m@     @Y@      $@      @      @      @              @      (@       @      ,@      &@      9@      @               @     �U@     `e@      @      &@     �Y@      7@     �n@     �J@     �j@     @X@      $@      @      J@      T@       @      .@     �\@      1@     �Z@     �K@     @_@     �V@      &@      @      ;@      I@      @      @     �U@      (@     �V@      A@      Y@      K@       @              @      ,@                      4@       @      <@      @      9@      @       @      @      8@      B@      @      @     �P@      $@      O@      ;@     �R@     �I@      @      �?      9@      >@      @       @      <@      @      0@      5@      9@     �B@      @      �?      "@      *@              @      0@      @      @      .@      0@      =@      @              0@      1@      @      @      (@      �?      $@      @      "@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJބ�/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�
(,;O@�	           ��@       	                    �?�P�z�@h           *�@                          �;@ǁj�b/@�           �@                           �?h�XmW@k           ��@������������������������       ���m��@	           �y@������������������������       ��哃(�@b            @c@                            �?L?(/��@-            �R@������������������������       ��8Ni�@             *@������������������������       ��w*�T@&            �N@
                           �?B'�9	@�           L�@                          �7@Ĺt�p@            y@������������������������       ��\!v�8@�            pq@������������������������       ��D��g@Q            @^@                           �?ܶ_Ӝ	@�           �@������������������������       �ƕAw�*
@�           І@������������������������       �o�rI/�@	           �z@                          �7@�Ok�:f@A           К@                           @�i�@@B           ��@                          �4@����@O           ��@������������������������       ��d!�� @�           ��@������������������������       ��[�K@�            0p@                           @Z�P�@�            �x@������������������������       ���ʖ�1@~             j@������������������������       ���d��i@u            �g@                            �?����y@�            @y@                           �?��l�@             i@������������������������       �C� �'@"             L@������������������������       �l�ᛮ�@]             b@                          �:@��X��E@�            `i@������������������������       ��=�@L            �_@������������������������       ���9��@4             S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     ��@      6@     �N@     �}@      Q@     Ȏ@     @n@     ��@     �w@      <@      2@     �h@     s@      .@     �C@     �s@      H@     �w@     �i@      x@     �p@      ;@       @     �L@     �R@      �?      @     �S@      @     �d@      @@     @c@      P@      @             �I@     @Q@      �?      �?     �P@      @      d@      7@      b@      F@      @              E@      L@      �?             �J@      @     @Y@      4@      Y@      A@      @              "@      *@              �?      ,@      �?     �M@      @      F@      $@               @      @      @               @      &@              @      "@      $@      4@       @       @      @      @                                                               @       @               @      @               @      &@              @      "@      $@      2@              0@     `a@     �l@      ,@      B@     �m@     �E@     @j@     �e@      m@     @i@      6@       @      1@      N@      �?       @      R@      @      Q@     �@@     �Q@      O@      @      �?      ,@      H@               @      H@       @     �H@      6@      L@      =@       @      �?      @      (@      �?              8@       @      3@      &@      ,@     �@@      �?      ,@     �^@     @e@      *@      <@     �d@     �C@     �a@     �a@     @d@     �a@      3@      ,@     �W@     �X@      *@      3@     �Y@      ;@     @P@     �Y@     �V@      U@      2@              ;@     �Q@              "@     �O@      (@     @S@      C@     �Q@      L@      �?      @      U@      p@      @      6@     �c@      4@     �@     �B@     Py@     �\@      �?             �M@     @j@      @      ,@     �X@      *@     ��@      7@     r@      P@      �?             �A@     �a@      �?      �?      H@      $@     �y@      ,@      j@      F@                      9@     �V@              �?      5@      @     �s@      &@     �c@      ?@                      $@     �H@      �?              ;@      @      Y@      @      I@      *@                      8@     �Q@      @      *@      I@      @     @^@      "@     @T@      4@      �?              2@     �@@              @      9@      �?     �S@      @     �B@      @                      @     �B@      @       @      9@       @     �E@      @      F@      ,@      �?      @      9@      H@      �?       @      M@      @     �R@      ,@      ]@      I@                      *@      A@              @      1@      @      B@      @      L@     �@@                       @      "@                       @      @      .@      �?      1@      @                      &@      9@              @      .@      �?      5@      @     �C@      ;@              @      (@      ,@      �?      @     �D@       @      C@      $@      N@      1@              @       @      @                      5@              6@      @      G@      *@                      @      @      �?      @      4@       @      0@      @      ,@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��|��b@�	           ��@       	                    �?�<���@n           *�@                           �?�˴s�@           0�@                          �<@^��$�@�            �r@������������������������       ��?wi@�            `q@������������������������       ���D��@             9@                           @&�X�`	@[           ��@������������������������       ��(�J0%	@1            @������������������������       �p�3�.�@*            @Q@
                           �?��+��@O           ��@                           �?�ߒ`d�@�            u@������������������������       �`j-�d@�            `o@������������������������       ���ݟu�@7            �U@                           �?y���-�	@x           ��@������������������������       ��P����	@�           ؆@������������������������       ��T5�+@�            0p@                           �?E����*@4           К@                          �4@F�� @l           0�@                            �?��z��3�?�            �u@������������������������       �-���t�?1            �T@������������������������       ��<�����?�            �p@                          �6@�l�@�            �l@������������������������       �<�x�,v@9            �W@������������������������       �ø�^Z7@P             a@                           �?����b@�           ��@                          �3@p=�݅n@\           ��@������������������������       ��mH�6�@�            @j@������������������������       �Sb���@�            �u@                           �?���nv@l           �@������������������������       �܃��@            �H@������������������������       ���Ȑ`�@R           `�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     0t@     Ѐ@      >@     �E@     P{@     �S@      �@     `n@     h�@     v@     �A@      7@      n@      s@      5@      A@      s@      L@     pw@     @h@     Pw@     `n@      <@      $@     @X@      `@      (@       @      `@      5@     �d@     @Q@     @_@      Y@      @              ?@      C@       @      �?     �A@      @     �U@      0@     @P@      :@                      >@      @@       @      �?      A@      @     @U@      *@      O@      0@                      �?      @                      �?              �?      @      @      $@              $@     �P@     �V@      $@      @     @W@      2@     �S@     �J@      N@     �R@      @      "@     �J@     �V@      @      @      T@      .@      S@      B@      I@      Q@      @      �?      *@      �?      @              *@      @       @      1@      $@      @              *@     �a@      f@      "@      :@      f@     �A@     `j@     @_@      o@     �a@      5@             �F@     �I@               @      B@             �R@      .@     @T@      ;@      @             �C@      E@               @      @@             �H@      ,@     �H@      6@       @              @      "@                      @              :@      �?      @@      @      @      *@     �X@     �_@      "@      8@     �a@     �A@      a@     �[@     �d@      ]@      0@      *@     @P@     �T@       @      4@     �\@      >@      S@      U@     @_@     @X@      0@             �@@      F@      �?      @      9@      @      N@      :@      E@      3@              �?     �T@      m@      "@      "@     �`@      6@     h�@     �H@     �{@     �[@      @              ,@     @T@              �?      ?@      @     0r@      (@     @_@      5@                      "@     �B@              �?      &@             @i@      @      S@      &@                              @                       @              K@              3@      @                      "@      A@              �?      "@             �b@      @     �L@      @                      @      F@                      4@      @     @V@       @     �H@      $@                      �?      4@                      (@      @      F@      �?      "@      @                      @      8@                       @       @     �F@      @      D@      @              �?     @Q@     �b@      "@       @     �Y@      0@     �t@     �B@     �s@     @V@      @      �?      ;@     �R@      @      @     �O@      @     @b@      3@     �d@     �G@      @               @      8@              �?      1@             @U@      @     �N@      "@              �?      3@      I@      @      @      G@      @     �N@      ,@     @Z@      C@      @              E@     @S@      @      @     �C@      &@      g@      2@     �b@      E@      �?                       @               @      @      @      (@       @      (@                              E@     @Q@      @       @      B@      @     �e@      $@      a@      E@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�:dehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?O�l@�o@�	           ��@       	                    �?�����	@�           @�@                          �6@��`��
@+           �}@                           �?�x���@�            r@������������������������       ���W��@I            �^@������������������������       � C#n�@n            �d@                           �?���<O@t             g@������������������������       ���R!�@,             R@������������������������       ����le�@H             \@
                          �:@�55c>"
@�           ܑ@                           @��UQ>
@)            �@������������������������       ��/��	@           `�@������������������������       ����Qt@             4@                           @Hl�5�	@�            �n@������������������������       ���I�ڃ	@&            �O@������������������������       ��ۥ5K�@r             g@                           @�`}�@�           �@                          �5@B�8��@i           X�@                          �1@|]j��L@�            �t@������������������������       ��.�A@9            �U@������������������������       �O�U�@�            �n@                            �?�zk� �@�             p@������������������������       �Ф!��7@*            �Q@������������������������       ������@l            @g@                           �?�[�j1@=           ��@                            �?}`�v�W@j           ��@������������������������       �X��e@�            �s@������������������������       ����/$�?�            0p@                           @�ۉW @�           ȑ@������������������������       ���al��@           ��@������������������������       ��Ao�S1@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        =@     0s@     �@      @@      N@     �y@     �T@     �@      i@      �@     �w@     �A@      <@     �g@     �m@      5@     �C@     �j@      H@     @l@     �^@     Pp@     @i@      :@      �?      K@     �S@      @      (@      G@      �?      W@      6@     @Z@     �L@       @              ?@     �I@      @      @      3@              Q@      *@     �R@      :@                      @      ;@                      @              ?@      @      G@      @                      8@      8@      @      @      .@             �B@      "@      =@      6@              �?      7@      ;@              "@      ;@      �?      8@      "@      >@      ?@       @      �?      *@      &@                       @              0@      �?      *@       @      �?              $@      0@              "@      3@      �?       @       @      1@      7@      �?      ;@     �`@      d@      2@      ;@      e@     �G@     �`@     @Y@     �c@      b@      8@      1@     �Z@      `@      .@      6@     ``@     �B@      ]@     �R@      a@     @W@      3@      (@     @Z@      `@      .@      6@      `@      B@     �\@     @R@      a@     �V@      ,@      @       @                               @      �?       @      �?               @      @      $@      <@     �@@      @      @     �B@      $@      2@      ;@      3@      J@      @      @       @       @      �?      �?      @      @               @      $@      &@      @      @      4@      9@       @      @      A@      @      2@      3@      "@     �D@      �?      �?     �]@     0s@      &@      5@     `h@      A@     �@     �S@     ��@     `f@      "@             �G@     @T@       @      $@      Q@      @     @b@      C@      `@     �L@       @              *@     �C@       @      @      A@      @     @Z@      1@     �T@      =@                      �?      .@                      @             �A@      @      3@      @                      (@      8@       @      @      ;@      @     �Q@      &@     �O@      9@                      A@      E@              @      A@      @     �D@      5@     �G@      <@       @               @      2@              @      @      �?      .@      @      $@      @       @              :@      8@              �?      <@       @      :@      2@     �B@      8@              �?     �Q@     @l@      "@      &@     �_@      ;@     x�@      D@     �{@     �^@      @              2@     �Q@      @      @      <@      @      q@      @     `a@      7@      �?               @     �C@      @       @      7@      @     �`@      �?      S@      5@                      $@      @@              �?      @             `a@      @     �O@       @      �?      �?     �J@     `c@      @       @     �X@      6@     �u@     �@@     0s@     �X@      @      �?      C@      ]@      �?       @      R@      *@     pq@      2@     �k@     �K@       @              .@     �C@      @      @      ;@      "@     �Q@      .@      U@      F@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJk�{zhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?v�XNVl@�	           ��@       	                    �?k�'V��@           ��@                           �?M����@>           ��@                          �1@�m��@w            @g@������������������������       ����+lY�?            �A@������������������������       ���~�{@c            �b@                          �5@��+A�@�            �u@������������������������       ���ws��@d            @f@������������������������       ��:�+�@c            �d@
                            @��¥�'@�           ؆@                            �?��^�s�@~           ��@������������������������       ��ǽ�� @r            �e@������������������������       �7�\+�@           {@                           �?6G���?T            @_@������������������������       �\���JT�?+             Q@������������������������       ��]�ٽ.�?)            �L@                          �1@ɾ{�=S@�           ��@                           @�V����@�            pv@                           @���Nx@!            �J@������������������������       �ߥf��@             9@������������������������       ��r�Vu��?             <@                          �0@��#O�@�             s@������������������������       ����@A             Y@������������������������       �C9���@�            �i@                           �?ݢ���@�           �@                           �?ّ��*	@q            �e@������������������������       �M��q!@"            �K@������������������������       �,ȥ¶	@O             ^@                           @<�MN�@O           ��@������������������������       ���h�6@�           ��@������������������������       �r���!�	@�            `q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     `t@     P�@     �C@     �G@     `|@     �U@     P�@      n@     ؇@     �v@      =@              W@     �e@      @      @     �]@      ,@     |@      H@     �p@     @V@      @             �N@     �U@       @      @     @R@      @     @`@      ?@      S@     �L@      @              6@      8@                      <@             �N@      @      >@      0@       @                      �?                      @              7@              @      �?                      6@      7@                      5@              C@      @      ;@      .@       @             �C@     �O@       @      @     �F@      @     @Q@      <@      G@     �D@      �?              3@      9@              @      3@      @     �H@      $@      >@      4@                      4@      C@       @      @      :@              4@      2@      0@      5@      �?              ?@     @U@      �?             �F@      &@     �s@      1@     �g@      @@      �?              <@      U@      �?              =@      &@     `o@      0@     @c@      ?@      �?               @      4@      �?               @      @     @T@              G@      "@      �?              :@      P@                      5@      @     @e@      0@      [@      6@                      @      �?                      0@              Q@      �?     �A@      �?                      @      �?                      (@             �@@              2@      �?                                                      @             �A@      �?      1@                      (@     @m@     �w@      B@      D@      u@      R@     H�@      h@      @      q@      9@              4@      L@               @      5@       @     @`@      *@     �T@     �@@                      @      @                      �?              8@      @      @      @                      @      �?                      �?               @      @      �?      @                      @       @                                      0@              @      �?                      *@     �J@               @      4@       @     �Z@      @      S@      <@                      @      >@              �?      @             �@@       @      ,@      &@                      "@      7@              �?      .@       @     @R@      @      O@      1@              (@     �j@     `t@      B@      C@     �s@     �Q@     pz@     `f@      z@     �m@      9@      @      7@      <@              &@      :@       @      $@      1@      ?@      1@      �?      �?       @      5@                      "@               @       @      $@      @      �?       @      5@      @              &@      1@       @       @      .@      5@      $@              "@     �g@     �r@      B@      ;@     r@      O@     �y@     @d@     x@     �k@      8@      @     �c@     �o@      >@      :@     `o@      H@     �w@     �_@     0v@     �g@      .@      @     �A@     �E@      @      �?      C@      ,@     �@@     �A@      >@      ?@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�p�e@�	           ��@       	                    �?�I��+	@&           �@                           �?(�x E�@/           `}@                          �9@�︐uj@x            �f@������������������������       �c�V��T@a             b@������������������������       �A �W}d@            �B@                            �?�D��u�@�            r@������������������������       ����Q�@:            �W@������������������������       �Z��3�@}            `h@
                           @(���	@�           ��@                           @��e�0n	@�           ��@������������������������       ���`�^	@�           ��@������������������������       �ĭ;�x�@�            Pq@                           �?Q���Ȟ@W            �`@������������������������       ��KD �@            �F@������������������������       �5_�m"0	@:            @V@                           �?�/��@�           ��@                            �?�z�f�@�           ��@                           �?_nV��@z            �g@������������������������       �ְ�!��??            �X@������������������������       �@��|n@;            @V@                          �5@��첇@X           ��@������������������������       ���@^A @�            @w@������������������������       ���7�,�@p             e@                           @�W�-8@�           ��@                          �1@<ݺ�M@�            �@������������������������       ���&H@D            �Y@������������������������       �z�܈�@q           Ё@                           �?4'D ��@           p�@������������������������       �O�ժ�K@           �z@������������������������       �����1@           Pz@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �p@     ��@      A@     �I@     �~@      T@     ��@     `j@     x�@     �v@     �A@      8@     �c@     �p@      5@      >@     @q@     �F@     @l@      a@     `p@     `i@      8@      �?     �E@     �P@      @      @     @Q@      @      [@      6@     �X@     �H@      �?      �?      2@      8@                      :@             �H@       @     �F@      0@                      &@      *@                      8@              F@       @      D@      $@              �?      @      &@                       @              @              @      @                      9@      E@      @      @     �E@      @     �M@      4@      K@     �@@      �?              "@      9@              �?      "@       @      2@      @      2@       @                      0@      1@      @      @      A@      @     �D@      0@      B@      9@      �?      7@     @\@     �h@      2@      :@     �i@      D@     �]@     �\@     `d@     @c@      7@      (@     �Y@     `e@      2@      9@     �f@      C@     @[@     @W@     �c@     �a@      ,@      (@     @S@     @]@      1@      *@     �b@      B@     �R@     �N@     �^@     @Y@      @              :@      K@      �?      (@     �@@       @     �A@      @@      B@     �C@      @      &@      $@      ;@              �?      :@       @      "@      5@      @      ,@      "@      �?      @      "@                      (@      �?              (@      �?      @      �?      $@      @      2@              �?      ,@      �?      "@      "@      @      $@       @              \@     �t@      *@      5@     �j@     �A@     ��@     �R@     H�@     �c@      &@              <@     @W@       @      �?      L@      @      u@      (@     `d@      @@       @              �?      5@       @      �?      1@             @T@       @      I@      &@       @                      @              �?      ,@              G@              9@      @                      �?      ,@       @              @             �A@       @      9@      @       @              ;@      R@                     �C@      @     �o@      $@     @\@      5@                      ,@     �J@                      8@       @     �h@      @     �P@      *@                      *@      3@                      .@      �?     �M@      @      G@       @                      U@     �m@      &@      4@     �c@      @@     0z@     �O@     `v@     @_@      "@             �A@     �^@      @       @      U@      :@      d@      F@     �^@     �M@      @               @      .@                      @             �F@      *@      0@      @                     �@@     �Z@      @       @      T@      :@      ]@      ?@     �Z@      J@      @             �H@      ]@       @      (@     �R@      @      p@      3@     `m@     �P@       @              :@     �K@      @       @      D@      �?     �`@      @     @^@      @@       @              7@     �N@      @      @     �A@      @      _@      0@     �\@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ#�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��é�S@�	           ��@       	                   �;@W`c�p6	@�           d�@                           �?1�l^��@=           �@                            @Vڣ�N@           �y@������������������������       �M�� *�@�            �o@������������������������       �ʥG4@d             d@                           @J�vd�m	@8           @�@������������������������       �����F	@,           ��@������������������������       �̴]E=@             3@
                           @���g�	@�            @q@                           �?:ס	�	@�             o@������������������������       ��J�Tq@-            @T@������������������������       ��p#�s@g            �d@                            �? .�ߵ@             <@������������������������       ��m�O�@
             .@������������������������       ��hfs���?             *@                           �?ad*�\@�           �@                           @P°�<@�           ��@                            �?��D��r@^           Ѐ@������������������������       �6#�;� @f            �c@������������������������       ���0�{@�            �w@                           �?�p$��m@�            �j@������������������������       ��Ip��V@L             ]@������������������������       ����@7            �X@                            �?�@�            �@                           @�V/,@�            v@������������������������       ������@I             [@������������������������       �&�F�c�@�            �n@                          �4@�5o>@�           |�@������������������������       �F��)@g           Ё@������������������������       �hnl@�           (�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     ��@     �@@      G@      }@     �Q@      �@     �k@     ��@     �u@     �B@      5@     �f@      k@      9@      ;@      p@     �A@     `n@     �_@      p@     �i@      =@      &@     @b@     �f@      1@      6@     `l@      9@     @k@      [@     �l@     �a@      9@              G@      N@       @      @     �H@      �?      Y@      ;@     �W@      :@      @              A@      >@      �?             �@@      �?     �O@      *@     �O@      (@      @              (@      >@      �?      @      0@             �B@      ,@      @@      ,@              &@      Y@     @^@      .@      2@     @f@      8@     �]@     @T@     �`@     �\@      6@       @     �W@      ^@      .@      2@      f@      8@     �]@     @S@     �`@     �\@      3@      @      @      �?                       @                      @                      @      $@      A@      B@       @      @      ?@      $@      9@      3@      =@     @P@      @      @     �@@     �@@       @      @      ;@       @      1@      ,@      <@     @P@      @      @      $@      "@      �?              ,@              .@      @      &@      *@               @      7@      8@      @      @      *@       @       @      &@      1@      J@      @      @      �?      @                      @       @       @      @      �?              �?       @              �?                      �?       @       @      @      �?              �?      �?      �?       @                      @              @                                              a@     Pt@       @      3@      j@     �A@     h�@      X@     x�@      b@       @              >@     �V@       @      @     �F@      @      u@      7@      g@      <@      �?              9@     �L@              �?     �@@      @     �o@      *@     �`@      .@                      @      7@              �?      @      �?     �R@             �C@       @                      4@      A@                      ;@      @     @f@      *@      X@      @                      @     �@@       @      @      (@             �U@      $@     �H@      *@      �?              @      3@              @      @              J@       @      5@      $@                       @      ,@       @              @              A@       @      <@      @      �?             �Z@     `m@      @      .@     `d@      <@     �y@     @R@     pw@     @]@      @              =@     �M@      �?       @      9@      @      \@      *@     @S@      <@                      @      :@               @      &@      @      :@      @      *@      (@                      7@     �@@      �?              ,@       @     �U@      @      P@      0@                     @S@      f@      @      *@     @a@      5@     �r@      N@     �r@     @V@      @              6@      [@       @      @     �H@       @     �f@      6@     �a@     �B@                     �K@      Q@      @       @     @V@      3@     �]@      C@     `c@      J@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJv��ehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@]1Ӂp@�	           ��@       	                    �?��o/�@t           6�@                           �?��r1@�           `�@                            �?�H��@           �z@������������������������       �A�Ͽz� @C            �]@������������������������       �,�����@�            `s@                           @1�')B�@�            �w@������������������������       �}�	�@�            `j@������������������������       ���ʠ��?p            �e@
                           @ܠ�b�@x           ��@                          �1@aq�,@�           ؆@������������������������       �E�h5�@q            �e@������������������������       ��+�:M@k           h�@                           @�] ��@�           ��@������������������������       �S;%n��@           �z@������������������������       ��Tԯ�@�            @m@                           �?(�?�i�@D           ��@                           �?�.枣@/           @                          �<@eW��k�@�            �o@������������������������       �n�}@}            �i@������������������������       ���(4�@#            �I@                           @�Y��@�            @n@������������������������       �&���/�@T             b@������������������������       ��\^�,@;            @X@                           @0q�*�m	@           ��@                          �9@>s�W�	@�           ȇ@������������������������       ���wu'	@           0y@������������������������       � C�Rp	@�            `v@                           �?�=�>ۭ@)           @|@������������������������       ������@�            `i@������������������������       �/9W���@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     X�@      >@     �O@      |@     �U@     p�@      m@     0�@     pv@      9@      @     @`@     �r@       @      >@     �k@      >@     `�@     �U@     0@     �d@      $@              L@     �X@              @     @P@      @     `u@      9@     �f@      >@      @              <@     �C@              @      D@      @     �i@      4@     @S@       @      @                      &@               @      &@      �?     �L@      @      >@      @                      <@      <@               @      =@      @     �b@      0@     �G@      @      @              <@      N@              �?      9@              a@      @     �Z@      6@                      7@     �A@              �?      2@              L@       @     �L@      3@                      @      9@                      @              T@      @     �H@      @              @     �R@     �h@       @      9@     �c@      :@     `w@     �N@     �s@      a@      @      @     �I@     �\@      @      ,@      _@      .@     @`@      H@     @_@      W@      @      @      (@      A@      �?      @      5@      �?      I@      "@      :@      *@              @     �C@     @T@      @      $@     �Y@      ,@      T@     �C@     �X@     �S@      @              7@      U@      @      &@      A@      &@     �n@      *@     �g@      F@       @              2@      I@      �?      @      <@      @     `d@      @     @`@      6@                      @      A@       @       @      @      @     @T@       @     �N@      6@       @      (@     �f@     p@      6@     �@@     `l@     �L@      r@     `b@     0q@      h@      .@       @      D@     �U@      @      @      L@      *@     @_@      >@     �X@     �A@      @       @      =@      J@       @      @      C@      �?      C@      2@      G@      8@      �?       @      8@      F@       @      �?      =@      �?      C@      .@      B@      &@      �?              @       @              @      "@                      @      $@      *@                      &@      A@       @              2@      (@     �U@      (@     �J@      &@       @              &@      .@                      @      $@     �L@      &@      <@      @       @                      3@       @              *@       @      >@      �?      9@      @              $@     �a@     `e@      2@      =@     `e@      F@     �d@     @]@      f@     �c@      (@      @      X@     �\@      (@      6@     @]@     �B@      O@     @W@     �S@     �\@      "@             �H@     �Q@      @      1@      Q@      2@     �E@      F@      G@      D@       @      @     �G@      F@      @      @     �H@      3@      3@     �H@      @@     �R@      @      @      G@     �L@      @      @      K@      @     �Y@      8@     �X@      F@      @      @      7@      @@              @      =@       @      D@      "@     �D@      .@      @              7@      9@      @      �?      9@      @     �O@      .@     �L@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ[�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�ml��`@�	           ��@       	                    �?փi�P�@n           ^�@                          �<@>Q���@�           @�@                            �?_�5$@n            �@������������������������       �A�O�A@�            �s@������������������������       ����"�@�            Pr@                            �?s��vr@/             R@������������������������       ��Hַ� @
             1@������������������������       �d����I@%            �K@
                           �?[� ��	@�           �@                          �2@�t+��	@�           ��@������������������������       �`v��@x             h@������������������������       �<��x>
@U           P�@                           �?��Vw��@           �y@������������������������       ���h @             A@������������������������       ���H�g)@�            �w@                           @	Ӹ ��@K           h�@                           �?�P��@�           t�@                           �?���W7��?�            �w@������������������������       ���!@��?�            `j@������������������������       ������f�?k            �d@                           @���qK@�           �@������������������������       �e��j��@�            `q@������������������������       �����vr@W           h�@                           @��C�
�@U           �@                           @���}�@�            �u@������������������������       �6qZ�@�            pp@������������������������       �%ŕuN�@9            �U@                           �?�0�n�~@h            �c@������������������������       ���ext@)             O@������������������������       �9���@?            @X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     0t@     P�@      9@     �N@     �y@     �T@     ȏ@      m@     Ȉ@     �v@      8@      8@      m@     �t@      2@      G@     �q@     @Q@      x@     @g@      w@      p@      5@              O@     �[@      �?      *@     �R@      @     �d@      E@     �a@      N@      @              N@     �W@      �?      @      P@      @      d@      B@     �`@     �D@      @             �A@      G@      �?      @      ;@       @     @S@      4@     @T@      2@      @              9@     �H@               @     �B@      @      U@      0@      K@      7@                       @      0@              @      $@              @      @      @      3@      �?              �?       @                       @                              �?      @      �?              �?       @              @       @              @      @      @      .@              8@     @e@     �k@      1@     �@@     �j@      P@     @k@      b@     @l@     �h@      1@      8@     �`@      c@      0@      9@     �c@      I@     ``@     @[@     �d@     �b@      1@              3@      3@              �?      9@      @     �A@      7@      F@      5@      �?      8@     �\@     �`@      0@      8@     ``@      G@      X@     �U@      ^@     @`@      0@              B@     �P@      �?       @      L@      ,@     �U@     �A@      O@     �G@                      @      @              @      @      �?              �?      @      @                      >@     �O@      �?       @     �H@      *@     �U@      A@     �M@     �D@              @     �V@     �k@      @      .@      `@      ,@     ȃ@      G@     �z@     �Y@      @      @      N@     �b@       @       @      U@      "@     �~@      7@     �q@     �O@      @              &@      D@                      0@      @     �k@      �?     �S@      @                      @      5@                      $@      �?      `@      �?      F@      �?                      @      3@                      @      @     @W@             �A@      @              @     �H@     �[@       @       @      Q@      @      q@      6@      j@     �L@      @      @      9@     �G@      �?      �?      >@      @     �R@      (@     �I@      ;@      �?              8@     �O@      �?      �?      C@             �h@      $@     �c@      >@       @              ?@     @R@      @      *@      F@      @     @a@      7@     @a@     �C@                      8@      I@      @       @      6@      @      \@      1@      W@      3@                      *@     �B@       @       @      0@      @      V@      0@     �P@      ,@                      &@      *@      �?              @              8@      �?      :@      @                      @      7@       @      @      6@       @      :@      @      G@      4@                      �?       @               @      "@      �?      @      @      1@      .@                      @      .@       @      @      *@      �?      4@      @      =@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@Oe3 �f@�	           ��@       	                    @���M])@y           d�@                           �?Ź�:V@6           ��@                           �?Ք7�{�@�            �r@������������������������       �U�2�?@W            `a@������������������������       ��U�-�@e            �c@                          �1@$+��d@z           ��@������������������������       ��z7@k            �e@������������������������       �7\xU��@           pz@
                          �1@����@C           ،@                           @g*7��?�            v@������������������������       �|����?;            �W@������������������������       �!^�I� @�             p@                           �?LC�G�@f           Ё@������������������������       ���v��?w            @f@������������������������       ������@�            �x@                          �;@l�l���@8           `�@                           �?�s�Rf@)           �@                          �9@^Jh��L@)           �}@������������������������       ��:ހ;@�            x@������������������������       �]���7@:             V@                           @���#Z�@            ��@������������������������       ���o� �	@�           x�@������������������������       �{'���,@0           �}@                           �?2�/6}	@           �z@                            �?Ⱦݽa�	@�            @p@������������������������       �T}=��;	@)            @P@������������������������       ��P��K	@w            `h@                           @?".cvV@o            �d@������������������������       ���cl�@2            @Q@������������������������       �몵G@=            @X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �r@      �@      ;@     �N@     �|@      V@     ��@     �i@     (�@      v@      =@      @     �U@     �o@      "@      ,@     �f@      0@     ��@     �T@     �x@     �a@      @      @     �J@     @_@      @       @     �_@      0@      k@     @Q@     �e@      V@      @              (@      F@              �?      >@       @     �X@      ,@      S@      2@                      @      3@                      3@       @      I@       @      8@      ,@                      "@      9@              �?      &@             �H@      @      J@      @              @     �D@     @T@      @      @     @X@      ,@     �]@     �K@     @X@     �Q@      @       @      *@     �@@      �?      �?      1@              H@      (@      @@      0@              @      <@      H@      @      @      T@      ,@     �Q@     �E@     @P@      K@      @              A@      `@      @      @     �K@             py@      *@     �k@     �J@                      @      D@              @      1@             `g@      @     �T@      0@                      �?      (@                      �?              P@       @      &@      @                      @      <@              @      0@             �^@      �?      R@      (@                      >@      V@      @      @      C@             �k@      $@     �a@     �B@                      "@      6@                      @             �V@      @      E@      @                      5@     �P@      @      @      A@              `@      @     �X@      ?@              4@     �j@     pt@      2@     �G@     pq@      R@      x@     �^@     �w@     `j@      6@       @     �e@     q@      ,@      <@     �j@     �F@     �u@      X@     �s@     �`@      6@             �G@     �U@       @       @     �D@       @     @b@      ,@      Y@      8@      @              G@     �O@       @       @      @@      @     �_@      ,@     �R@      1@      @              �?      7@                      "@      @      3@              9@      @               @     @_@     `g@      (@      :@     `e@     �B@     �i@     �T@      k@     @[@      3@      @      X@     �^@       @      8@      ^@      ;@     �S@      N@     �V@     �Q@      .@      �?      =@      P@      @       @     �I@      $@     �_@      6@     �_@      C@      @      (@      E@      K@      @      3@     �P@      ;@     �A@      ;@     �N@     �S@              (@      <@     �@@       @      .@      =@      3@      (@      8@      =@     �L@              @      @      *@              �?      @       @      @      @      @      "@               @      6@      4@       @      ,@      7@      &@      @      2@      6@      H@                      ,@      5@       @      @      C@       @      7@      @      @@      5@                      �?      ,@       @      @      $@      @      @      @      .@      $@                      *@      @                      <@      @      0@              1@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJa�+JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @s:��5)@�	           ��@       	                    �?�}63Ӧ@�           h�@                            �?�Z	�d�@           ��@                           �?yo�-'�@3            ~@������������������������       �����@a            �b@������������������������       ��J��u#@�            �t@                           @�Վ"0	@�           $�@������������������������       ��x�\c�@�           ��@������������������������       ��Ox�5@6            �V@
                           �?oj]�9@o           H�@                            @�;G��;@v            �g@������������������������       ��L���~@Z            `b@������������������������       ������?            �D@                           �?�D���@�            �x@������������������������       ���cu&@             B@������������������������       ��ƁA\@�            �v@                           @I]�@F           T�@                           @r�S)�T@-           ��@                           �?7����@$           ��@������������������������       ��X����?�            �w@������������������������       �<$���{@5           @}@                           @���#�O@	           �y@������������������������       �F?��$�@�            �o@������������������������       ���jD�E@`            �c@                            @��_O��@           �z@                           @F�ӂ@�            Pv@������������������������       ���P2��@�            u@������������������������       �8���N�@             4@                           @�ڪ�h�@)            @Q@������������������������       ��y��@             2@������������������������       �V���%�@            �I@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      s@     h�@      5@     �L@     �{@     �S@     ��@     �i@     `�@     �v@      ?@      .@      k@     Pt@      ,@     �F@     �t@     �P@     `y@     �e@     w@     �n@      7@      .@     �d@     �n@      *@      @@     �o@      J@     �n@     @^@     0q@     �i@      6@      �?      H@     �N@      �?       @     @U@      @      S@     �E@     �X@      G@      $@              ,@      =@               @      1@      �?     �A@      @     �A@      &@      @      �?      A@      @@      �?      @      Q@      @     �D@     �C@     �O@     �A@      @      ,@     �]@     �f@      (@      8@     �d@     �G@      e@     �S@      f@     �c@      (@      @      ]@     @e@      (@      8@     �b@      F@     �c@     �P@     �e@     �a@      "@       @      @      *@                      2@      @      $@      (@      @      1@      @             �H@     @T@      �?      *@     �S@      .@      d@     �I@     �W@     �D@      �?              3@      *@                      3@      @     @S@      @      F@      @      �?              1@      (@                      $@      @     �L@      @     �B@      @      �?               @      �?                      "@              4@              @       @                      >@      Q@      �?      *@     �M@      (@      U@      F@      I@      B@                      @      @               @      @              @      @      @      @                      :@     @P@      �?      @      K@      (@     @T@     �B@     �G@     �@@              @      V@      m@      @      (@     �\@      (@     @�@     �A@     �{@     �\@       @      @      I@     �e@      @      (@     @T@       @     `~@      >@      u@     �Q@       @      @      =@     �Z@      �?      @      K@      @     pv@      *@     �l@     �E@                      &@     �G@                      $@              g@      @     �Z@      .@              @      2@     �M@      �?      @      F@      @     �e@      @     @_@      <@                      5@     �P@      @      @      ;@      @     �_@      1@     �Z@      <@       @              "@     �G@       @      @      3@      @     �Q@      *@     �P@      0@       @              (@      3@      @      @       @             �L@      @      D@      (@                      C@      N@      �?              A@      @     @`@      @     @Z@     �E@      @              >@     �L@                      >@       @      Z@      @      W@     �@@      @              8@     �L@                      :@             �Y@      @     @V@      >@      @              @                              @       @      �?      �?      @      @                       @      @      �?              @       @      :@              *@      $@       @              @                              �?              @               @      �?       @              �?      @      �?              @       @      5@              &@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ކhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@ 3�5@�	           ��@       	                    �? W�L5S@W           �@                          �1@��C*�@�           ��@                          �0@���� @�            �n@������������������������       ��oy @:            �U@������������������������       �F�t�[<�?k             d@                          �4@|cjN@E           �@������������������������       �">å��@�             y@������������������������       �Q�<c�@H             Z@
                          �1@?���c@m           �@                           @h�I6�@�             v@������������������������       �{�D=��@k            `f@������������������������       � ��&�?n            �e@                           @M.���@�           ��@������������������������       �1���=@Z           ��@������������������������       �` \3~C@:            �@                           �?�%6�@Y           X�@                            �?��G�	�	@&           0�@                           �?y��O:�	@�            @q@������������������������       �ퟒj�@8             U@������������������������       ��G��[�	@z             h@                           �?Bfh���	@t           ��@������������������������       ��Z�K	�@y            �j@������������������������       �\����	@�            �w@                           @L:cR��@3           ��@                            @�X�@           X�@������������������������       �d�F��@�           X�@������������������������       �6)~24@w             h@                            �?(ٙ��.@            �B@������������������������       ����L&@             1@������������������������       �Pu�x�{@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      r@     ��@      =@      K@     �|@      U@     �@      i@     p�@     `w@      ;@      @      `@     �t@      @      3@     �h@      =@     �@     �R@     �}@     �f@       @              F@     �W@      �?       @     �E@      @     �t@      ,@      d@     �J@       @               @      :@               @      7@             �`@      �?     �C@      &@       @                      (@                      3@             �B@              ,@      @                       @      ,@               @      @             �X@      �?      9@      @       @              B@     @Q@      �?              4@      @      i@      *@     @^@      E@                      =@      J@                      3@       @     �c@       @     �W@      C@                      @      1@      �?              �?       @     �D@      @      :@      @              @     @U@     �m@      @      1@      c@      9@     @w@      N@     �s@     �_@      @              5@      P@       @       @      &@      @     �`@      &@     �S@      >@                      1@     �B@       @              @      @     �H@      &@      >@      7@                      @      ;@               @      @             �T@              H@      @              @      P@     �e@      @      .@     �a@      6@      n@     �H@     �m@     @X@      @      @     �F@     �W@      �?       @      X@      2@     @S@      E@     �W@     �K@      @              3@      T@      @      @      G@      @     `d@      @     �a@      E@       @      *@      d@     @m@      6@     �A@     pp@     �K@     t@     �_@     0s@     @h@      3@      (@     �X@     �`@      2@      4@     �a@     �A@      V@     �S@     �[@     @]@      ,@      @      @@      ?@      @      @     �L@       @     �C@      >@     �@@      9@      @              @       @      �?              7@      �?      .@      @      @      0@       @      @      9@      7@      @      @      A@      @      8@      9@      ;@      "@      @       @     �P@      Z@      *@      *@     �U@      ;@     �H@      H@     �S@      W@      "@       @      6@      A@       @      @      @@      @      <@      @      >@      C@      @      @     �F@     �Q@      &@      @      K@      4@      5@     �D@      H@      K@      @      �?      O@     �X@      @      .@      ^@      4@      m@      H@     �h@     @S@      @      �?     �I@      X@      @      .@      \@      3@     �l@      C@     @h@     @S@      @      �?     �D@      U@      @      &@      S@      3@      f@      >@     @c@     �I@      @              $@      (@      �?      @      B@             �K@       @      D@      :@                      &@      @                       @      �?       @      $@       @                              @      �?                       @      �?              @       @                              @       @                      @               @      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ�^>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�-�U@�	           ��@       	                    �?f8I�t�@�           x�@                          �<@���ZP�@�           8�@                          �5@�O���0@|           ��@������������������������       ����j�@�            �u@������������������������       �0�\z�G@�            �k@                          @@@�	�^u@2             T@������������������������       �g�� �@)            �P@������������������������       ��bN�� @	             ,@
                          �4@�{R�d	@�           Ԙ@                           �?L����b@~           ��@������������������������       ��""�*6@�            �j@������������������������       �����^	@�            �z@                           �?��4��	@X           ȍ@������������������������       ��~��/
@�           ��@������������������������       ����@�             m@                           �?E�5�&�@            4�@                            @����@j           ��@                          �>@�a٪˼@,           `}@������������������������       �rPY�[4@%           �|@������������������������       ��;N�@             *@                          �3@���<��?>            �V@������������������������       ���S����?$             K@������������������������       ��vs��?             B@                          �7@���D:�@�           t�@                           @aW�8�}@           X�@������������������������       ���[g@n            �e@������������������������       ��B�@��@�           ��@                           @@\�8��@�             s@������������������������       ��R�z�<@�            �q@������������������������       �d��B�@	             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     Ȁ@      ;@     �K@      |@     �U@     ȏ@     �l@     ��@     @w@      >@      .@      j@     Pt@      7@      F@     u@      O@     �w@     �g@     �v@     �p@      <@             �P@     @V@       @      @      V@      @     �d@      A@     @_@      N@      @             �K@     �S@       @      @     �R@      @      d@      :@     �]@      C@      @              3@     �C@       @      @     �D@      @      \@      2@     �S@      9@       @              B@     �C@               @     �@@      �?      H@       @      D@      *@      @              &@      &@               @      ,@              @       @      @      6@      �?              "@      "@              �?       @              @       @      @      6@      �?               @       @              �?      @                              @                      .@     �a@     �m@      5@     �B@      o@      L@     �j@     @c@     �m@     �i@      6@      @      F@     �R@      "@      1@      Z@      &@     @_@     �H@      [@     �U@      @       @      0@     �C@      @       @     �C@      @     �A@      2@      7@      <@               @      <@      B@      @      .@     @P@      @     �V@      ?@     @U@      M@      @      &@     �X@      d@      (@      4@      b@     �F@      V@     @Z@     @`@      ^@      2@      &@     �R@     �_@      (@      2@     �Y@     �@@     �O@     �R@     �W@      W@      2@              7@     �A@               @      E@      (@      9@      >@     �A@      <@               @     �W@     �j@      @      &@     @\@      8@      �@     �D@     �z@     �Z@       @              =@      N@               @      9@      @     �q@      (@     �_@      1@      �?              ;@     �L@              �?      8@      @     @l@      &@     @Y@      1@      �?              ;@      L@              �?      7@      @      l@      "@     @Y@      (@      �?                      �?                      �?       @       @       @              @                       @      @              �?      �?             �L@      �?      9@                               @                                              A@              2@                                      @              �?      �?              7@      �?      @                       @     �P@      c@      @      "@      V@      3@     Pv@      =@     �r@     @V@      �?             �B@     �]@      @      @      G@      *@     pr@      &@     �k@      N@      �?              @      @@                      &@      "@     �N@      @     �B@      ,@      �?              @@     �U@      @      @     �A@      @     @m@      @      g@      G@               @      =@      A@      �?      @      E@      @      O@      2@      T@      =@               @      9@      @@      �?      @     �B@       @      N@      ,@      T@      =@                      @       @                      @      @       @      @                        �t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ!�(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�R?)�(@�	           ��@       	                    @�̓�-@@@           ��@                           �?V����@�           ��@                          �<@��
U��@           @z@������������������������       ��gB#Z�@�            0x@������������������������       ���;l�]@            �@@                          �4@XG�w�@�           ��@������������������������       �Lu��@�            �s@������������������������       ����a��	@           `|@
                            �?�(kgb�@U           �@                          �5@�Xb�*�@�            x@������������������������       ���/Ě��?�            �n@������������������������       �ƶ̾v@X            �a@                           @(�@q~T@]            �@������������������������       �1.����@M            @[@������������������������       �_��v�f@           0{@                           �?�:����@y           �@                          �;@��+ۄ�@r           �@                          �3@*��Z.@M           H�@������������������������       �RDJCv�@�             o@������������������������       ��&�J?�@�             q@                          �=@�jo7�@%             M@������������������������       �M�2��T@             >@������������������������       �� ڭ@             <@                           @�a5��@           �@                           �?�U`l"	@           H�@������������������������       ��f��	@W           @�@������������������������       �e6>��/@�            r@                           �?�ō�!�@�            �y@������������������������       �rN[S݇@
             2@������������������������       ��|P>�4@�            �x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �q@     ��@      =@      M@     0z@     �S@     h�@     �i@     `�@     @v@      ;@      3@     �b@     �q@      &@     �@@     �h@      H@     P�@      `@     �}@     �h@      0@      3@      Z@     �d@      "@      >@     �`@      @@     �j@     �Z@     �m@     �^@      .@       @      A@     @P@      �?      $@      H@      (@     �T@      H@     �P@      C@      @       @      ?@     �M@      �?      $@      F@      "@     �T@      E@     �P@      ;@      @              @      @                      @      @              @              &@              &@     �Q@     �X@       @      4@     �U@      4@     @`@     �M@     @e@      U@       @              ;@     �B@      @      �?     �A@      @     �S@      3@      R@      @@      @      &@     �E@      O@      @      3@      J@      1@      J@      D@     �X@      J@      @              F@     �^@       @      @      P@      0@     Pu@      6@     �m@     �R@      �?              4@     �D@                      :@      @     �e@      (@     @T@      ;@                      @      8@                      (@             `a@      @      J@      @                      ,@      1@                      ,@      @     �A@      @      =@      5@                      8@     @T@       @      @      C@      (@     �d@      $@     �c@      H@      �?              @      .@              �?      @      (@     �@@      �?      8@      (@      �?              4@     �P@       @       @      @@             �`@      "@     �`@      B@              @      a@     �q@      2@      9@     �k@      ?@      @     @S@     u@     �c@      &@              D@     �S@      �?      @     �M@       @      m@      ,@     @[@     �B@      �?             �@@     �N@      �?      @     �G@       @     `l@      &@     @Y@     �@@      �?               @      3@              @      5@      �?     @^@      @      K@      0@      �?              9@      E@      �?      �?      :@      �?     �Z@      @     �G@      1@                      @      1@               @      (@              @      @       @      @                      @      .@                       @               @      �?      @      �?                       @       @               @      $@              @       @      @      @              @     @X@     `i@      1@      3@      d@      =@     �p@     �O@     �l@     �^@      $@      @      V@     `a@      ,@      .@     @]@      :@      `@      L@      _@     �U@      $@      @      N@     �T@      *@      (@     @V@      2@     @P@     �B@     �Q@     �L@      $@      �?      <@      L@      �?      @      <@       @     �O@      3@     �J@      =@                      "@      P@      @      @      F@      @      a@      @      Z@      B@                       @      @               @      �?      @       @      �?       @                              @     �M@      @       @     �E@             �`@      @     �Y@      B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����~}@�	           ��@       	                    �?��f��@�           ��@                           �?�;�дI@�           �@                           �?�+�t��@0           `|@������������������������       �>'f�@~            �g@������������������������       �e�5cgw@�            �p@                           �?L�⍝@r            �f@������������������������       ��*)�@@5            @U@������������������������       �;p[� @=            �X@
                          �5@��&��	@�           @�@                          �0@��ג)�@�           ��@������������������������       ���A��u@             K@������������������������       ��ۣq��@�            �@                           �?��e�x�	@           Њ@������������������������       �U�=}%@.            @U@������������������������       ��l�76�	@�           (�@                           @(NOo4@           �@                           @l�c� @�           �@                          �7@�
}�@�           ��@������������������������       �֏���@p           x�@������������������������       ��;ւ:2@Z            �a@                          �5@Bw3�� @           �y@������������������������       ������?�            r@������������������������       ��;A��P@U            �_@                          �6@wK���@N           �@                           @�[Ś�7@�            0u@������������������������       �_1��=_@�             t@������������������������       ��{�V�@
             1@                           @˗�g @u            �e@������������������������       ���F�r*@A            �X@������������������������       � �<q k@4            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     pu@     Ѐ@     �@@      Q@     �{@     �S@      �@     �k@     ؉@     v@      A@      *@     �o@     Pt@      8@      L@     �s@     �O@     �v@     �f@     Py@     �l@      :@      �?     @Q@     �R@      @      @      V@      @     �a@      B@     @d@     �I@      @      �?      L@     @P@      @       @     @Q@      �?     �U@      ?@     �W@      D@      @      �?      .@      :@                      ?@             �E@       @      H@      0@       @             �D@     �C@      @       @      C@      �?      F@      7@     �G@      8@       @              *@      $@              �?      3@       @     �K@      @     �P@      &@                      @      @              �?      .@      �?      >@      @      3@      @                      @      @                      @      �?      9@      �?      H@      @              (@      g@     @o@      5@     �J@     �l@      N@     @k@      b@     `n@      f@      6@      "@     �I@     @]@      @      :@      ]@      .@      a@      O@     �a@     �Q@       @              @      4@              �?      @              $@              @      "@              "@      G@     @X@      @      9@     �[@      .@     �_@      O@      a@     �N@       @      @     �`@     �`@      ,@      ;@     �\@     �F@     @T@     �T@     �Y@     �Z@      ,@       @      4@      "@               @      .@      �?      �?      @       @      (@       @      �?     �\@      _@      ,@      3@      Y@      F@      T@     �R@     �W@     �W@      (@      �?     @V@     �j@      "@      (@     @^@      0@     ��@      D@     `z@     @_@       @      �?     �M@      b@       @      @     �Q@       @     �|@      6@     r@     @T@      @      �?      F@      X@       @      �?      G@       @     �p@      4@     �f@      N@      @              @@     �T@       @             �@@      @      n@      ,@     �a@      B@      @      �?      (@      ,@              �?      *@      @      <@      @     �C@      8@                      .@      H@              @      9@              h@       @     �Z@      5@                       @      >@              @      @             �b@             �T@      (@                      @      2@                      4@             �F@       @      9@      "@                      >@     @Q@      @      @      I@       @     �a@      2@     �`@      F@      @              2@     �G@       @      @     �@@       @     @[@       @      X@      6@      @              1@     �F@       @      @      =@       @     @[@       @     �W@      3@                      �?       @              �?      @                               @      @      @              (@      6@      @      @      1@      @      A@      0@     �B@      6@                       @      1@      @      @      @       @      5@      *@      6@      "@                      $@      @       @              $@      @      *@      @      .@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�l��y@�	           ��@       	                    �?A�-�	@S           ��@                           �?נD��	@�           d�@                          �;@�sf1�@0           P~@������������������������       ������@           0y@������������������������       ��
���@.            �T@                           �?��2�;�	@�           Б@������������������������       � <y�U�@           �y@������������������������       ��6$�_
@�           Ȇ@
                          �3@+�RBs@^           (�@                           �?b G��@{            �h@������������������������       �{��Z� @'            �N@������������������������       �!��6oF@T             a@                          �<@�d/@�            �u@������������������������       �����@�            �s@������������������������       ������@            �A@                           @Z	~��@L           ,�@                          �2@�zp-@�           ̒@                           @u�G,ώ�?           �{@������������������������       ��¼cs��?�             v@������������������������       ����<o�?;             V@                           @"��j��@�           ȇ@������������������������       ���>'-@/           �}@������������������������       �����@�             r@                           �?*pP��@S           ��@                          �6@P����@�             l@������������������������       �N�6@]            @c@������������������������       �����g�@,            �Q@                           �?��$�5@�            �s@������������������������       �R ��5@^            �b@������������������������       �v��q��@l            @d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �r@     ��@     �A@     �K@     �|@     �V@     l�@     �l@      �@     @w@      <@      8@      k@     �s@      :@      C@     s@      Q@     �w@     @h@     �t@      o@      :@      8@     �f@      l@      9@      >@     �m@      I@     �n@     �a@     �l@     `j@      8@      �?      K@     @S@       @      "@     @P@      @     �Y@      @@      U@      I@       @              G@      P@       @      @     �I@      @      X@      =@     �R@      ?@       @      �?       @      *@              @      ,@      @      @      @      "@      3@              7@      `@     �b@      7@      5@     �e@     �E@     �a@     �[@     `b@      d@      6@       @      4@      N@      @      @     @P@      *@     �Q@     �D@      O@     �N@      @      5@      [@      V@      0@      .@     �Z@      >@     �Q@     @Q@     @U@      Y@      3@             �A@     �V@      �?       @      Q@      2@     �`@      J@     �Y@     �B@       @              "@      A@                      ,@             �P@      0@     �G@      &@                      @      @                       @              0@      �?      <@      @                      @      >@                      (@             �I@      .@      3@      @                      :@     �L@      �?       @      K@      2@      Q@      B@     �K@      :@       @              6@     �H@      �?      @     �G@      0@     �P@      ;@      K@      8@       @              @       @              �?      @       @      �?      "@      �?       @               @     �T@     �j@      "@      1@     `c@      7@      �@      A@     py@      _@       @       @      L@     �a@      @      @     @X@      0@     �@      3@     `q@      R@      �?              &@     �D@      �?              2@             �m@             �^@      &@                      &@     �@@      �?              2@             @g@              Y@      @                               @                                      J@              6@      @               @     �F@     �Y@       @      @     �S@      0@     q@      3@     �c@     �N@      �?       @      A@      K@       @       @     �M@      0@      b@      .@     �W@     �H@      �?              &@      H@              @      4@              `@      @      O@      (@                      :@     @Q@      @      (@      M@      @      d@      .@      `@      J@      �?              @      9@      �?      @      .@      �?     �X@      @      L@      ,@      �?              @      1@              @       @             @T@      @      =@      @      �?                       @      �?              @      �?      1@      �?      ;@       @                      7@      F@      @      @     �E@      @     �O@      $@     @R@      C@                      "@      7@      @      @      6@      @     �@@      @      >@      2@                      ,@      5@       @      �?      5@      @      >@      @     �E@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @iU���@�	           ��@       	                    @qT�,@�           ��@                          �8@>���@W           �@                           �?����G@`           ��@������������������������       �-Z��@�            �s@������������������������       �5[u��	@�           ��@                           �?��#Rx	@�            y@������������������������       �-�θ��@_            `c@������������������������       ���"^�	@�            �n@
                          �7@��%�S@|           D�@                            �?0He��9@�           ��@������������������������       ��LG�jd @�            pr@������������������������       �p����@�           ��@                            �?�_h	�%@�            0u@������������������������       ��o�ׄ@}            @i@������������������������       ���Wv��@V             a@                           �?����H@�           ؑ@                          �:@n䌟F	@�           (�@                          �6@G�&��k@p           ��@������������������������       ��	��\1@�            �y@������������������������       �.����F@s            �c@                           @׶)�t
@M             a@������������������������       �.�<��D
@8            @V@������������������������       �����@             H@                           �?@�P
�@           {@                          �3@����?T            �a@������������������������       �b����?-             R@������������������������       ��iM�� @'             Q@                           @r+mD6@�            Pr@������������������������       �;A�h�@J            �Z@������������������������       �F�:y�@v            `g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     Ps@     ��@      A@      G@     p|@      Y@      �@     �i@     ��@      x@     �A@      (@     �h@      x@      2@      >@     0r@      S@     `�@      b@     �@     �p@      9@      (@     �`@     �g@      @      3@     `f@     �N@     �k@     �[@      n@      c@      5@      @      X@     @`@      @      1@     �]@     �A@     @g@      P@      h@      V@      @              >@      D@      �?              B@      @     �Y@      "@     �R@      3@      @      @     �P@     �V@      @      1@     �T@      @@      U@     �K@     �]@     @Q@      @      @      C@      M@      �?       @      N@      :@     �A@      G@     �H@     @P@      ,@       @      $@      ?@      �?      �?      5@      @      ,@      7@      *@      =@      @      @      <@      ;@              �?     �C@      3@      5@      7@      B@      B@      &@             @P@     �h@      &@      &@      \@      .@     �~@      A@      w@     �\@      @             �G@     @c@      &@      @     �P@      $@     @{@      0@     �p@     @Q@       @              "@     �@@      @              (@              c@       @     �P@      *@                      C@     @^@      @      @      K@      $@     �q@      ,@      i@      L@       @              2@      E@              @      G@      @     �M@      2@      Y@     �F@       @              @      3@              @      6@      @      D@      $@     �Q@      :@                      &@      7@              �?      8@      �?      3@       @      =@      3@       @      0@     �[@      b@      0@      0@     �d@      8@      o@     �N@     �j@     @]@      $@      0@     �T@      X@      (@      *@      `@      2@      W@     �D@     @]@     �T@      $@      @      N@     @T@       @      @      [@      *@     �T@     �A@     �Z@      N@       @      @      H@      I@      @      @      M@       @     �Q@      :@     �U@     �I@      @              (@      ?@      @       @      I@      @      *@      "@      3@      "@      @      (@      7@      .@      @      @      5@      @      "@      @      &@      6@       @      @      &@      *@      @      �?      2@      @      @      @      $@       @       @      @      (@       @              @      @               @      @      �?      ,@                      ;@     �H@      @      @     �A@      @     �c@      4@     �X@     �A@                      &@      @                      &@             �R@      @      ?@      @                      @      �?                                     �D@              5@      @                      @       @                      &@              A@      @      $@      �?                      0@      G@      @      @      8@      @     @T@      0@     �P@      >@                      $@      9@       @      �?      @       @      7@      (@      ,@      *@                      @      5@       @       @      4@      @      M@      @     �J@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?@6�ԛ4@�	           ��@       	                    �?��"b�@           d�@                          �<@�y�2��@;           �~@                          �9@�5J��@           �{@������������������������       �
ߖ�3h@�            0x@������������������������       ��d�a@$            �J@                           �?�'!x��@%            �J@������������������������       �>�u��@             :@������������������������       �އ��F�@             ;@
                            �?16� �{@�           `�@                          �7@��Ѐ @z             g@������������������������       ��[�����?e            `c@������������������������       �HVc�6 @             =@                            @����@j           ��@������������������������       ��YB��@           �{@������������������������       �Ɨ0����?V            �^@                           @ �ԁ@�           �@                          �2@�5�3	@�           �@                           �?��n�@�            t@������������������������       ���V��/@|            @j@������������������������       ��^�� �@C            �[@                           �?�/�ێ	@            �@������������������������       �NK6�N�@�            0t@������������������������       ��6s	f�	@L           �@                           �?�2�(G�@�           ��@                           @����mB@I           `@������������������������       �=���}@�            `t@������������������������       �tj���@s             f@                           @dJ��N@m           ȁ@������������������������       ��$�m?@�            0x@������������������������       �fť��@q            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     ؁@      :@     �D@     �|@      W@     h�@     �i@     �@     w@      <@      �?     �T@     �h@      @      &@     �Y@      .@     pz@      D@     �q@     �R@      @      �?     �H@      W@       @      @     �L@      @     �X@      :@     @[@      G@      @      �?     �E@     �T@       @      @     �H@      @     �W@      7@     �Y@      ?@      @             �C@     �P@       @      @      C@       @     �U@      4@     �W@      >@      @      �?      @      .@                      &@      �?      "@      @       @      �?                      @      $@               @       @              @      @      @      .@                              "@              �?      @              �?      �?      @       @                      @      �?              �?      @               @       @      @      @                      A@     �Z@      �?      @      G@      (@     Pt@      ,@      f@      <@      �?                      6@      �?      �?      @      @     �V@      �?      H@      $@                              6@      �?      �?      @      �?     �T@             �A@      @                                                      �?       @       @      �?      *@      @                      A@      U@              @     �C@      "@     @m@      *@      `@      2@      �?              ?@     �S@               @      ?@      "@     @e@      (@      W@      ,@      �?              @      @              �?       @              P@      �?     �B@      @              2@     @j@     Pw@      7@      >@     @v@     @S@     0�@     �d@     (�@     pr@      8@      1@     �b@     �l@      4@      6@     @n@     @P@     �l@     �a@     p@      j@      4@      �?      9@      A@       @             �K@      @     �S@      <@     �N@      @@      �?      �?      7@      7@       @             �D@       @      C@      0@     �C@      8@      �?               @      &@                      ,@      �?     �D@      (@      6@       @              0@      _@     �h@      2@      6@     `g@      O@     �b@      \@     �h@      f@      3@      �?      .@      J@              @     �I@      "@      L@      :@      I@     �K@       @      .@     @[@      b@      2@      0@      a@     �J@     �W@     �U@     @b@     �^@      1@      �?     �N@     �a@      @       @     �\@      (@      t@      ;@     @r@     �U@      @      �?      8@     �S@       @      @     @Q@      @     `a@      *@     @`@      @@      @      �?      &@     �L@              @     �F@       @     @S@       @     @[@      3@                      *@      6@       @       @      8@       @      O@      &@      5@      *@      @             �B@      P@      �?      @     �F@       @     �f@      ,@     @d@      K@                      7@     �I@               @      9@      @     �`@      @     �\@      :@                      ,@      *@      �?      �?      4@      @      G@      @      H@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�w;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���;Ɔ@�	           ��@       	                   �<@~��V�"	@�           z�@                           �?��X���@�            �@                          �;@/��d)�@�           ��@������������������������       �	�焊O@z           8�@������������������������       ����@
             (@                           @�-�q�	@o           ԕ@������������������������       �Ⱦ.�q	@R           �@������������������������       �, ����@            �G@
                           @-@J}�b	@�            �n@                          �=@�rd��	@L            �_@������������������������       ��%����@             E@������������������������       � ���=
@1            @U@                           @ӵ�h�$@J            �]@������������������������       �|V/�o@>            �X@������������������������       ���'�,�@             3@                            �?>�Q�@<           0�@                          �5@� �K�7@�            @x@                          �4@hDw��v�?�             n@������������������������       �dI�6XA�?�            �j@������������������������       �*#S���?             ;@                          �8@d��8��@]            �b@������������������������       ����)�@/             S@������������������������       �*r��@.             R@                           @
�Oe'@@            �@                          �2@P� �y@?           ��@������������������������       ��2�a�!�?�            Pu@������������������������       ��A'�@k           8�@                            @�����@           �x@������������������������       ����F�.@�            �p@������������������������       ���s�!@Q             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     ��@      D@      M@     z@     �V@     `�@      l@     ��@     �u@      >@      8@     �m@     `t@      >@      E@     `r@     �Q@     v@      g@     �x@     �o@      :@      2@     �j@     �q@      :@      ?@     pp@      J@     �u@     @d@     Pw@     �h@      8@      @      O@     �T@      �?      @      R@      @     �d@      5@      a@     �E@                     �N@     @T@      �?      @     �Q@      @     @d@      5@      a@     �E@              @      �?       @                      �?      �?      @              �?                      .@      c@     �i@      9@      ;@     �g@      H@     �f@     �a@     �m@      c@      8@      &@     �a@     `i@      9@      ;@     @g@     �G@     `f@     �`@     @l@     �b@      3@      @      $@      �?                      @      �?       @      @      $@       @      @      @      8@     �C@      @      &@      ?@      3@      @      6@      8@      L@       @      @      2@      1@      @      $@      4@      @      @      $@      &@      8@      �?              (@      @       @      �?      �?              �?       @      @      .@              @      @      *@       @      "@      3@      @      @       @      @      "@      �?       @      @      6@              �?      &@      0@       @      (@      *@      @@      �?              @      4@              �?      "@      $@       @      "@      *@      =@               @               @                       @      @              @              @      �?      �?     �R@     @n@      $@      0@     �^@      4@     X�@     �D@     y@      W@      @              ,@      H@       @              3@      @     `f@       @     �T@      =@                      �?     �@@                       @              `@      @     �K@      &@                      �?      :@                      @              _@      @     �E@      $@                              @                       @              @              (@      �?                      *@      .@       @              &@      @      I@      @      <@      2@                      $@      "@       @               @      @      >@              @       @                      @      @                      @      �?      4@      @      8@      $@              �?     �N@     @h@       @      0@      Z@      ,@     �}@     �@@     �s@     �O@      @      �?      C@     ``@      �?      �?     �M@      $@     0w@      2@      l@     �A@       @              &@     �E@      �?              "@             �e@      @      V@      (@              �?      ;@      V@              �?      I@      $@     �h@      ,@      a@      7@       @              7@     �O@      @      .@     �F@      @     @Y@      .@     @W@      <@       @              1@     �G@      @      @     �A@      @      M@      *@      O@      1@       @              @      0@      �?       @      $@      �?     �E@       @      ?@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@R��6W@�	           ��@       	                   �1@\̐��@�           ��@                           �?~:�*~@�           ��@                          �0@̵�1D�?�            �n@������������������������       ����G��?1            �U@������������������������       �d��0��?k            �c@                            �?6K�3�@�             v@������������������������       �6�w�@7            @S@������������������������       ��Xd�0@�            Pq@
                           �?ﭓe�@           �|@                           @,`WW�@t             i@������������������������       �~�^��@@            @Z@������������������������       ��A��@4             X@                           �?�R���"@�            `p@������������������������       ��7��I@;            �V@������������������������       �.DiXS�@b            �e@                           �?��#�]1@           H�@                          �<@�N�9Cp@           ��@                            @t
Z*ɧ@�           ��@������������������������       �n�j�@K           �@������������������������       �*.�.��@�            @k@                          �>@��7P)�@6            �X@������������������������       �����]@              N@������������������������       �4��vn+@            �C@                          �<@�hZM�@           ��@                           @ik��@~           @�@������������������������       ��b�b�	@�           �@������������������������       ��5�,��@�           h�@                           @�B�	�	@�            �k@������������������������       �l?��	@m            �c@������������������������       �����z�@+             O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @q@     `�@      =@     �O@      {@     �Q@     Џ@     `l@     @�@     0w@     �C@             �J@     `c@      �?      &@     �U@      @     @y@     �C@     �l@      R@      @              7@     �U@              @     �D@      �?     p@      ,@     �`@     �A@      �?              @      @@              �?      *@             ``@      �?     �I@       @      �?                      .@                      @              E@      �?      4@      @                      @      1@              �?       @             @V@              ?@      @      �?              1@      K@              @      <@      �?     �_@      *@      U@      ;@                      �?      "@                      $@      �?      D@       @      $@      @                      0@     �F@              @      2@             �U@      &@     �R@      7@                      >@     @Q@      �?      @     �F@      @     `b@      9@     �W@     �B@      @              ,@      <@      �?              <@      �?     �P@      @     �F@      &@       @              &@      5@                      3@      �?      9@      @      1@      @       @              @      @      �?              "@             �D@              <@      @                      0@     �D@              @      1@      @     @T@      4@      I@      :@       @              @       @              @      *@      �?      *@      0@      .@      (@       @              &@     �@@              �?      @       @      Q@      @     �A@      ,@              5@     �k@     y@      <@      J@     �u@     �P@     0�@     �g@     �@     �r@      A@      �?      N@      ^@      @       @     �Q@       @      p@      =@     �h@     �P@      @      �?      L@     �Y@      @      @     �I@      @      o@      3@     �f@      G@      @      �?     �C@     �P@       @      @     �E@      @      f@      (@     @_@      <@      @              1@      B@      �?      @       @              R@      @      L@      2@                      @      1@              �?      3@      �?       @      $@      0@      5@       @               @      0@                      @              @      @      &@      ,@       @               @      �?              �?      ,@      �?      @      @      @      @              4@     `d@     �q@      9@      F@     `q@      M@     `v@     �c@     �w@      m@      =@      ,@     �a@     @o@      5@      C@      o@      F@     �u@     �`@     Pv@     �g@      ;@      (@     @Y@     �d@      *@     �@@     �e@     �A@     �`@     @Y@     �f@     @_@      5@       @     �C@     @U@       @      @     �R@      "@     �j@     �@@      f@     �O@      @      @      7@      ?@      @      @      >@      ,@      &@      9@      8@      F@       @      @      $@      3@       @      @      3@      ,@      @      9@      ,@      B@       @              *@      (@       @      �?      &@              @              $@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ0�rwhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @*��fV@�	           ��@       	                    �?���/��@m           V�@                           �?o����0	@�           ��@                          �<@Cڇ��S@�           ��@������������������������       �Ԏ�A�%@^           ��@������������������������       �^=�*@"             L@                           �?ɒ7�m	@a           P�@������������������������       �B��N@�            �q@������������������������       �^��y��	@�           ��@
                           �?��`2�@�           h�@                          �7@��1�{@�            �p@������������������������       �]���(�@u            �g@������������������������       �!s2�QI@3             T@                          �2@]���B@�            �u@������������������������       ��ӴAy@?            @X@������������������������       ��a� @*@�            �o@                           @V���Q@2           x�@                           @o
#��c@�           |�@                            �?7XZ��@�            �y@������������������������       ������@�            �m@������������������������       ���p�@i            �e@                           �?A��HW@�            �@������������������������       ��f�*'�?�             m@������������������������       �� &<�@_           ؀@                          �8@y����@B           �@                           �?��p@�g@�            px@������������������������       ���z�^@h            @e@������������������������       ���X���@�            �k@                           �?�]��wi@N             ^@������������������������       ���[�@             �I@������������������������       ��&!^@.            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     s@     p�@      D@      H@     `{@      U@     ��@     �h@     �@      x@      A@      .@     �j@     �s@      >@      ?@     �r@     �P@     �w@     �d@     `y@     �p@      <@      .@     �d@     �l@      <@      =@      l@      F@     �l@      \@     �q@     �j@      :@      @     �E@     @V@      @      &@     @Y@      &@      _@     �B@     @[@     �S@      .@      @      B@     �U@      @      &@      Y@      $@      ]@      A@     �Y@     �K@      .@              @      @       @              �?      �?       @      @      @      8@              &@     �^@     �a@      7@      2@      _@     �@@     @Z@     �R@     �e@     �`@      &@              <@     �J@      �?      @      =@      �?     �G@      5@     �O@      >@      �?      &@     �W@     �U@      6@      &@     �W@      @@      M@      K@     @[@     @Z@      $@              H@     @U@       @       @      S@      6@     @c@     �J@     @_@      J@       @              7@      <@      �?      �?      C@      ,@     �K@      :@     �M@      9@      �?              $@      7@      �?      �?      ?@      ,@     �D@      4@     �E@      @      �?              *@      @                      @              ,@      @      0@      3@                      9@     �L@      �?      �?      C@       @     �X@      ;@     �P@      ;@      �?               @       @                      @      �?     �G@      @      6@      @                      7@     �H@      �?      �?      A@      @      J@      4@      F@      5@      �?             �V@     �n@      $@      1@      a@      2@     ��@     �@@     pz@     �]@      @             �J@     �f@      @      @     @W@      ,@      |@      8@     �r@     �L@      @              4@      R@       @       @      <@      *@     @b@      (@     @V@      7@      @              ,@     �K@       @       @      &@      "@     �R@      @      F@      2@      @              @      1@                      1@      @      R@      @     �F@      @      �?             �@@      [@      �?      @     @P@      �?      s@      (@     @j@      A@      �?              @      :@                      @      �?     �a@      �?      I@      @                      =@     �T@      �?      @     �M@             �d@      &@      d@      =@      �?              C@      P@      @      (@      F@      @     `b@      "@      _@     �N@      �?              ?@      H@      @      @      :@      @     �`@      �?     �X@      B@      �?              &@      8@      �?      �?      @             �S@             �C@      &@      �?              4@      8@      @      @      6@      @     �L@      �?     �M@      9@                      @      0@       @      @      2@      �?      (@       @      :@      9@                      @      $@              @      @               @      @      "@      $@                      @      @       @      �?      .@      �?      @      @      1@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJS<=YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @UaɓV'@�	           ��@       	                    �?���)��@j           f�@                           �?nQ�Lr�@�           H�@                           �?��Y!WR@4           @������������������������       �@փ8@r            �g@������������������������       ���X@�            Ps@                          �<@$0�y�a@r             g@������������������������       ����0+@k            @e@������������������������       ��t}�c@             ,@
                          �5@-����7	@�           (�@                           �?�1�@�           ��@������������������������       �V��gb@B           x�@������������������������       ���Ld@�            @l@                           �?�fI��	@�           Ȉ@������������������������       ��dJ���@%             O@������������������������       �v�ӝ�	@�           ؆@                           �?N�+�@1           X�@                            �?�}<�� @j           8�@                           �?�@�=#d�?N            �`@������������������������       ��m34��?%            �M@������������������������       ��ފ$;q�?)            �R@                          �3@v�7�?� @            |@������������������������       ����L$�?�             m@������������������������       ��9����@�             k@                           @�ƛZ�@�           <�@                            @�m��@�           (�@������������������������       ������@�           �@������������������������       �9� �m @E             Z@                            �?��ÄY@�            �t@������������������������       �w��8ň@/            �U@������������������������       �cW4W��@�            `n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     ��@      >@      K@     �{@     �T@     ,�@     @j@     `�@     x@      8@      0@     `k@     `t@      1@     �F@     �s@     �O@     Pw@     �d@     x@     �q@      6@             �Q@      V@      @      $@      T@       @      c@      ?@     �c@      S@      @             �I@     �P@      @      $@     @Q@      @     �W@      8@     �Z@     @P@       @              *@      6@                      2@              K@      @     �J@      6@                      C@     �F@      @      $@     �I@      @      D@      2@     �J@     �E@       @              4@      5@                      &@      @     �M@      @     �I@      &@      �?              4@      2@                      &@      @      M@       @      I@       @                              @                                      �?      @      �?      @      �?      0@     �b@     �m@      *@     �A@     `m@     �K@     �k@     �`@     �l@     �i@      3@      @     �I@     �\@      @      (@     �[@      6@      a@     �K@     �`@     @Z@      @      @      E@      S@      @       @     �U@      0@     �R@     �A@     �W@     �T@      @              "@     �C@              @      8@      @      O@      4@      D@      6@              *@     @X@     �^@      "@      7@     @_@     �@@      U@      T@     @W@     �X@      ,@      @      $@      3@               @       @                      @      @      @      @      $@     �U@      Z@      "@      5@     @]@     �@@      U@     �R@     �U@     �W@      &@      �?      Q@     �i@      *@      "@      `@      4@     ��@      F@     �z@     @Z@       @              ,@     �R@       @              @@      @     `q@       @     �b@      1@                              1@       @               @      @     @R@              ;@       @                              @                       @      @      @@              0@       @                              *@       @              @      �?     �D@              &@                              ,@      M@                      8@      @     �i@       @     �^@      .@                      @      2@                      .@             �]@      @     �O@      "@                      "@      D@                      "@      @     �U@      @      N@      @              �?      K@     ``@      &@      "@     @X@      *@      x@      B@     Pq@      V@       @      �?      @@     @W@      @      @     @Q@      @     �r@      3@      g@     �L@       @      �?      >@     @V@      @      @      J@      @     �p@      3@     `b@      J@      �?               @      @                      1@             �B@              C@      @      �?              6@      C@       @       @      <@      "@     �T@      1@      W@      ?@                      @      @              �?      @      �?      ?@      @      ;@      @                      0@     �@@       @      �?      6@       @      J@      *@     @P@      9@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ2�rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?C�7S@�	           ��@       	                    @����c@           P�@                           �?!��4';@�           h�@                            �?O[_ּ@9           �~@������������������������       �:�����@X            @b@������������������������       �a�;��1@�            �u@                          �;@⊽ct�@l            �c@������������������������       �:�4�%@_            @a@������������������������       ��恃�@             5@
                           @WZV�� @o           8�@                          �9@�,q��?�            �r@������������������������       ��Q��D�?�            �o@������������������������       �&� LH@            �H@                           @�m��S�@�            �q@������������������������       ��C�ףG�?3            �U@������������������������       ���ZȶQ@z            `h@                          �3@�Ð�I@�           �@                           �?f!_�@2           h�@                            @��}��
@+            @Q@������������������������       �UD/<��@             H@������������������������       ��a��@             5@                          �1@���`�@           @�@������������������������       �1�c@�            Pu@������������������������       �	�J�|@.           0@                          �:@ .�x�@P           ��@                           @��؆��@E            �@������������������������       �]�Tzm@           ��@������������������������       �%�*�K@&           P}@                          �;@�gS�_�	@            z@������������������������       ����\h@H             [@������������������������       ���K�z�	@�            @s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     ��@     �A@     �M@     �|@     �R@     ��@     �k@     �@     v@     �@@      �?     �T@     �d@      @       @      \@       @     �{@      C@     Pr@     @R@      @      �?     @P@     @X@      @      @      V@      �?     �c@      =@     �b@      J@       @      �?     �I@     @U@      @      @     @Q@      �?     �Y@      9@      Z@      F@      �?      �?      "@      >@                      7@              >@      @     �B@      &@                      E@     �K@      @      @      G@      �?      R@      4@     �P@     �@@      �?              ,@      (@              �?      3@             �K@      @     �F@       @      �?              (@       @              �?      &@             �J@       @     �E@       @                       @      @                       @               @       @       @              �?              1@     �Q@      �?      �?      8@      @     �q@      "@      b@      5@       @              (@      @@                      @      @     �d@       @     @P@      $@                      (@      :@                      @      �?      b@       @      L@      @                              @                      �?      @      6@              "@      @                      @      C@      �?      �?      1@             @^@      @     �S@      &@       @              �?       @                      @              D@              <@      @                      @      >@      �?      �?      $@             @T@      @     �I@       @       @      0@     `i@     �x@      =@     �I@     �u@     �P@     ��@      g@     �@     �q@      =@      @     �C@     �\@       @      *@     �X@      $@     r@      K@     �g@      V@       @      �?       @      "@              @      *@       @      ,@      @       @      "@                              @                      "@       @      ,@      @      @      @              �?       @      @              @      @                      @      �?       @              @     �B@     �Z@       @      "@     @U@       @     0q@     �G@     �f@     �S@       @       @      0@      I@      �?       @      1@      �?     �^@      ,@     �T@      @@              �?      5@      L@      @      @      Q@      @      c@     �@@     �X@     �G@       @      (@     �d@     �q@      5@      C@      o@     �L@     @q@     ``@     �s@      h@      ;@       @      `@      l@      .@      ;@      g@      E@     �k@     �W@     0p@      `@      6@       @     �T@     �^@      $@      3@      ]@     �A@     @d@     �F@      g@     �W@      $@             �G@     �Y@      @       @     @Q@      @     �N@     �H@     �R@     �A@      (@      $@     �A@     �L@      @      &@      P@      .@     �J@     �B@      N@     �O@      @      @      @      @      �?       @      1@              :@      *@      .@      3@      �?      @      <@     �J@      @      "@     �G@      .@      ;@      8@     �F@      F@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJKE=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��r�k@�	           ��@       	                   �5@_��>k	@�           �@                          �1@V����@�           ��@                           @�t�p�P@h            �e@������������������������       �U�j4@T             a@������������������������       �ɸ݋�@            �A@                           �?���H�D@m           X�@������������������������       �+{=Z2�@�            @n@������������������������       �^�q{�@�            �u@
                           �?7V>�k6
@           �@                          �<@̸�8�@�            �l@������������������������       ���L|@u             f@������������������������       ��j���Z@"             K@                          �6@=��y
@}           ��@������������������������       �h��}f
@C            �Y@������������������������       ���Q0
@:           P@                          �1@q��/;@�           �@                            �?D	ѵ[� @           }@                           �?Ml/ @�            `p@������������������������       �S�J���?E            @]@������������������������       �G�{j�� @X             b@                           @nX�o{ @z            `i@������������������������       ���1�� @f            `e@������������������������       �*T�Ja��?             @@                           @��2��@�           ��@                          �;@���כ@F           0@������������������������       �����b@'           P|@������������������������       �31Y��@             G@                          �6@ ���
@>           ,�@������������������������       �|.�.`;@           ��@������������������������       �E�6���@9           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     @s@     0�@      @@     �R@     p}@      T@     �@     `l@     ��@     pu@      =@      .@     `f@     @j@      6@     �E@     �m@     �G@     �l@      a@     �o@     �h@      7@      @     �Q@     �Z@       @      *@     �[@      2@     �a@     �I@     �b@      U@      @       @      .@      :@                      .@             �D@      @     �B@      ?@                      "@      4@                      "@             �C@      @      A@      5@               @      @      @                      @               @              @      $@              @      L@     @T@       @      *@     �W@      2@     �Y@      G@     �\@     �J@      @      �?      0@      G@              @      E@       @     �D@      5@     �H@      1@               @      D@     �A@       @      @     �J@      0@     �N@      9@     @P@      B@      @      $@      [@     �Y@      4@      >@      `@      =@     @U@     @U@      Z@     @\@      3@       @      8@      A@              "@      ?@       @      C@      ,@     �F@      >@       @       @      5@      <@              �?      8@       @     �B@      $@      C@      (@       @              @      @               @      @              �?      @      @      2@               @      U@     @Q@      4@      5@     �X@      ;@     �G@     �Q@     �M@     �T@      1@       @      *@      $@      @       @      @      @       @      0@      .@      *@              @     �Q@     �M@      .@      *@     �V@      5@     �C@     �K@      F@     �Q@      1@       @      `@     @s@      $@      @@      m@     �@@      �@     �V@     ��@     @b@      @              &@      O@              @      9@              n@      &@     �W@      0@      �?               @      B@              @      4@              a@      @     �J@      @                      �?      1@              @       @              Q@              4@                              �?      3@                      (@              Q@      @     �@@      @                      "@      :@                      @             @Z@      @      E@      "@      �?              "@      3@                      @             �V@      @      A@      "@      �?                      @                                      .@       @       @                       @     �]@     �n@      $@      =@     �i@     �@@     x�@      T@     0{@     @`@      @             �C@     �R@       @      $@      R@      ,@     @\@      E@      W@      C@      @             �@@     �P@       @      $@     �O@      ,@     �Z@     �B@      U@      C@                      @       @                      "@              @      @       @              @       @     �S@     �e@       @      3@     �`@      3@     �{@      C@     pu@      W@       @             �B@      \@      @      @     �S@      (@     �r@      ,@      i@     �K@       @       @      E@      N@      �?      *@      L@      @     �b@      8@     �a@     �B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJFr5OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?����hx@�	           ��@       	                    �?i�%�sF@           4�@                           �?��c�h@B           @�@                            �?)=Ͷ�X@�            �h@������������������������       �$`ƙ��@-            @Q@������������������������       ����4X�@S             `@                          �3@�$S$o	@�             t@������������������������       �p��u�@C            �^@������������������������       ���CH@             i@
                          �5@`B��@�           (�@                           @s���[� @I           @@������������������������       ��������?�            �w@������������������������       ���k_n@S             ^@                           @���D�@�             j@������������������������       ��)��V2@U            �^@������������������������       ���Չ�@7            �U@                            @�D	�u2@�           ��@                           !@�˺�@�           0�@                          �7@�$d/��@�           �@������������������������       �Zj2(�@F           D�@������������������������       ��/L	@u           H�@������������������������       �~�G��	@             2@                           @����	@�           ��@                           �?4�Po�	@e           @�@������������������������       ���Y�	@           @}@������������������������       �>=<�4@H             ]@                          �9@��d�]�@n             e@������������������������       �}���@W             `@������������������������       �
y�}7A@             D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �s@     ��@     �A@      I@     �z@     �V@     @�@      j@     Ȉ@      w@     �A@      �?      T@     �g@      @      *@     �\@      .@     �z@     �H@     @n@     @U@      @      �?      L@      X@      @      "@     @P@      @     @Y@      @@     @W@     �L@      �?      �?      4@     �B@                      1@             �E@      (@      I@      2@              �?      @      (@                      @              3@              4@      @                      .@      9@                      (@              8@      (@      >@      &@                      B@     �M@      @      "@      H@      @      M@      4@     �E@     �C@      �?              @      ,@              �?      8@      @      >@      @      4@      4@                      >@     �F@      @       @      8@       @      <@      0@      7@      3@      �?              8@     �W@      @      @     �H@      $@     �t@      1@     �b@      <@      @              3@     �Q@              @      ?@       @     Pp@      $@     �V@      &@       @              &@      M@               @      7@       @      j@      @     �O@      @                       @      (@               @       @             �J@      @      ;@      @       @              @      8@      @              2@       @     �P@      @     �M@      1@      �?              @      0@                      @       @      E@      @      ;@      "@      �?                       @      @              &@              9@              @@       @              1@     �m@     �y@      <@     �B@     �s@     �R@     ؀@      d@     8�@     �q@      ?@      "@     �e@     �q@      (@      4@     �j@     �J@     �y@     �^@     0z@     �g@      3@      "@     @e@     �q@      (@      4@     �j@      H@     �y@     �^@      z@     �g@      0@      @     �Y@     �k@      @      .@     �b@      8@     Pu@     �P@     Ps@     �\@      "@      @      Q@     �N@      @      @     �P@      8@     �Q@     �K@     @[@     �R@      @              @       @                      �?      @              �?      �?              @       @      P@     �^@      0@      1@     �X@      6@     �_@     �B@     �`@      X@      (@       @      L@      [@      (@      1@     �U@      5@      S@      B@     @S@     @S@      $@       @     �E@     �S@      "@      0@     @S@      2@     �I@      9@      Q@     @P@      $@              *@      >@      @      �?      "@      @      9@      &@      "@      (@                       @      .@      @              (@      �?     �I@      �?     �K@      3@       @              @      .@      �?              @      �?     �D@             �E@      &@       @              �?              @              @              $@      �?      (@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�h;%�\@�	           ��@       	                    �?�ad�|@           <�@                          �6@Mk�7�@           �|@                          �3@"��	�@�            �p@������������������������       �!r\��f@g            �d@������������������������       ��q�9�@?             Y@                            �?��[$�	@v            @h@������������������������       ��:q��@F             _@������������������������       ��6��@0            �Q@
                          �>@pi�'�W@�           (�@                            �?��BQG� @�           ��@������������������������       �b���?v            `i@������������������������       ��R_O%�@f           h�@������������������������       ��0~�Ά@
             *@                          �5@D��H&f@�           ��@                           @��C��@l           �@                          �1@M����@           ��@������������������������       �=^v�K[@�            �s@������������������������       ���Y:@O           (�@                           �?"3��@R            �`@������������������������       �f)��v@             H@������������������������       �����@5             U@                           @3~�+r	@3           ��@                           �?�%�O�
@            �@������������������������       ���L�	@�            �h@������������������������       �r���"
@�            �@                           @S�����@!           @{@������������������������       �^ wۧf@           Pz@������������������������       ���}�@	             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        5@     0q@     P�@      >@     �I@     �z@      Z@     Џ@     `j@     p�@     Pw@     �A@       @     @R@     @d@      @      @      Y@      &@     �|@      D@     �r@      R@      @       @      C@     �Q@       @      @      O@       @     �U@      9@     @]@     �F@      @              6@     �E@       @      �?      9@      �?     @Q@      ,@     �P@      3@       @              @      @@                      5@      �?     �F@      @      C@      .@                      0@      &@       @      �?      @              8@       @      <@      @       @       @      0@      ;@              @     �B@      �?      1@      &@     �I@      :@      @       @      &@      ,@              @      6@      �?      (@      @      ;@      8@      @              @      *@                      .@              @      @      8@       @                     �A@      W@      �?      �?      C@      "@     pw@      .@     `f@      ;@      �?              A@     �V@      �?      �?      A@       @     pw@      &@     `f@      9@      �?              �?      5@      �?              @       @      Z@             �N@      @                     �@@     �Q@              �?      ;@      @     �p@      &@     �]@      3@      �?              �?      �?                      @      �?              @               @              3@     @i@     �x@      ;@      G@     pt@     @W@     h�@     `e@     0�@     �r@      =@      @     �R@      j@      @      4@     �b@      F@     �v@     @P@     pt@     �`@      (@      @     �P@      h@      @      3@     �`@     �@@     �t@      L@     �s@      ]@      @       @      0@      E@              �?      3@              \@       @      U@      =@              @      I@     �b@      @      2@      ]@     �@@     @k@      H@     �l@     �U@      @      �?      "@      0@              �?      .@      &@      ?@      "@      ,@      2@      @      �?      @      @                      "@      @              @      @      @      @              @      *@              �?      @      @      ?@       @      "@      &@      @      *@     �_@     �f@      4@      :@      f@     �H@     �h@     �Z@     �g@     �d@      1@      (@     �X@     �_@      1@      2@      ]@     �D@     �U@     @W@      Y@      \@      .@      �?      (@      ;@      @      @      <@      @      ?@      0@      <@     �A@      @      &@     �U@      Y@      ,@      (@      V@     �B@     �K@     @S@      R@     @S@      $@      �?      <@      L@      @       @     �N@       @     �[@      *@     �V@     �K@       @      �?      5@      K@      �?       @     �M@       @     �[@      (@     �V@     �K@       @              @       @       @               @                      �?      �?                �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�8_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���n�/@�	           ��@       	                     �?5V����@           L�@                           �?��w��W@�           `�@                            �?� �ŌC@�            �s@������������������������       �	�R�@]            @a@������������������������       �,,��K@r            `f@                          �6@R��@�            �t@������������������������       ����#"�@�             k@������������������������       ��/�mF@F            �]@
                          �3@H��͛@o           8�@                            @p��G� @�             q@������������������������       �ڏ8I�?E            @]@������������������������       �"i��� @[            `c@                           @�D
*�@�            ps@������������������������       �ӳ���@}             h@������������������������       ����� @R            �]@                           @G`m�	@�           �@                           @E7-	@�           ��@                            �?���X�	@�           ��@������������������������       �I<e��@�            �w@������������������������       �u�!Q�@�             v@                          �4@�
W.+�@�           ��@������������������������       �=aK^�o@�             s@������������������������       ���3G�	@.           �}@                          �7@V�
��@�           �@                            �?߮�G��@           ��@������������������������       �Tw�͡@t            �g@������������������������       ��07�O�@�           ��@                           �? l���@�            ps@������������������������       ���hɹ!@T            �\@������������������������       �e���C�@s            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     8�@      1@      I@     @}@     @W@     �@     @j@     ��@      u@     �@@      �?     �X@     �d@      �?      @     �]@      $@     @{@     �F@     �q@     �O@      "@      �?      J@     �W@      �?      @      O@      @      j@      5@     �b@     �F@       @      �?      2@      F@               @      9@      @     �\@      ,@      P@      8@      @      �?      @      *@                      (@       @      M@      @     �@@      &@                      ,@      ?@               @      *@      @     �L@      $@      ?@      *@      @              A@      I@      �?      �?     �B@       @     �W@      @     @U@      5@      @              7@     �@@                      &@              R@       @      O@      *@                      &@      1@      �?      �?      :@       @      6@      @      7@       @      @             �G@     �Q@              @      L@      @     `l@      8@     �`@      2@      �?              "@      .@                      .@       @     @a@      (@     �Q@      "@      �?               @      @                      @       @     �P@      @      9@       @      �?              @      "@                      "@             �Q@      @      G@      @                      C@      L@              @     �D@      �?     @V@      (@     �N@      "@                     �@@      B@              @     �B@      �?      B@      (@      >@      @                      @      4@              �?      @             �J@              ?@      @              1@      k@      x@      0@     �E@     �u@     �T@     ��@     �d@     �@     0q@      8@      1@      c@     `n@       @      :@     `m@      Q@     �j@     �`@      l@      f@      5@      *@      Q@      ]@      @      0@      [@      D@      \@     �B@     �^@     �V@      @      @     �F@     �K@       @      *@     �E@      <@      J@      3@     �R@     �F@               @      7@     �N@      @      @     @P@      (@      N@      2@      H@     �F@      @      @      U@     �_@      @      $@     �_@      <@     @Y@     �X@     @Y@     �U@      .@              1@     �D@       @              P@      @      O@     �A@      F@      :@      "@      @     �P@     �U@      �?      $@     �O@      6@     �C@     �O@     �L@     �N@      @              P@     �a@       @      1@     �\@      .@     �w@      >@     �q@     �X@      @              C@     �^@      @      $@      Q@      &@     �t@      $@     @i@      H@      @              1@      <@                      0@       @     @S@      @     �B@      "@                      5@     �W@      @      $@      J@      "@     �o@      @     �d@     �C@      @              :@      5@      @      @     �G@      @      I@      4@     �T@      I@                      .@      0@               @      2@              .@      @      >@      *@                      &@      @      @      @      =@      @     �A@      ,@      J@     �B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�n�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?5㍊K@�	           ��@       	                   �;@��i�		@           h�@                          �9@x�����@d           ��@                           @v�^ԛ@           �@������������������������       ���_)��@9           ��@������������������������       ��x@b��	@�            0s@                            �?��u�@`            �c@������������������������       �Æ�9@#             M@������������������������       ���a�5@=            @Y@
                          @@@dx�K�@�            �n@                          �>@�_"��@�            �i@������������������������       ���::w@h            �d@������������������������       �.I����@             D@                           @q��A�j@            �D@������������������������       �p�%�4�@             :@������������������������       ��^">� @	             .@                           @Њ<�@�           ޡ@                            �?ǼA�h�@j           �@                           �?�(>�f@o            �f@������������������������       �Mݖ
�+@+             R@������������������������       �@m�fG@D            @[@                           �?7(�4@�            �x@������������������������       ������@I             ^@������������������������       �����e	@�            @q@                            �?�c1pR@*           ��@                          �4@XX[Z'@I           ��@������������������������       ��k�z@G           ��@������������������������       ��7���@           �y@                          �4@�E3:��@�           ��@������������������������       �'vq�;@�            `x@������������������������       �H*p��3@�            `w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      q@     `�@      <@     �R@     �|@     �R@     0�@      j@     `�@     �u@      >@      2@      d@     �o@      *@     �D@     0q@     �D@     �i@      `@     �p@     �h@      6@      (@      a@     �k@       @     �A@      n@      >@      h@      [@     @n@     �`@      5@      &@     ``@      h@      @     �A@     �j@      7@      f@     �T@      k@     @]@      .@      @      X@      `@      @      5@     �d@      *@     �b@      H@      g@     �V@      @      @     �A@     �O@      �?      ,@     �G@      $@      <@     �A@      @@      ;@      &@      �?      @      >@      �?              <@      @      0@      9@      9@      .@      @               @       @                      $@      @      @      .@      ,@               @      �?      @      6@      �?              2@      @      (@      $@      &@      .@      @      @      9@      ?@      @      @      A@      &@      ,@      4@      =@      P@      �?      @      6@      4@      @      @      =@      &@      *@      4@      3@      M@      �?      @      3@      3@      @      @      ;@      $@      "@      "@      .@     �F@                      @      �?                       @      �?      @      &@      @      *@      �?      @      @      &@       @              @              �?              $@      @              �?      @      @       @               @                              $@      @               @              @                      @              �?                      @               @     �[@     �t@      .@      A@     @g@     �@@     ��@     @T@     �@     �b@       @              A@      W@       @      *@      M@      .@      c@      H@      ]@     �F@       @              @      >@              @      5@      @     �G@      .@     �D@      &@       @                      "@                      2@              6@      @      1@      @                      @      5@              @      @      @      9@      (@      8@       @       @              =@      O@       @      $@     �B@      "@     @Z@     �@@     �R@      A@                      "@       @                      @              I@       @     �A@      @                      4@      K@       @      $@      ?@      "@     �K@      9@      D@      >@               @     @S@     `n@      *@      5@      `@      2@     ��@     �@@     �z@     @Z@      @             �F@     �a@      @      &@      P@      (@     �u@      8@     �l@     @Q@                      5@     �M@      @      @      7@             �m@       @     �`@      D@                      8@     �T@              @     �D@      (@     @[@      0@     @X@      =@               @      @@     �Y@      "@      $@      P@      @     Pr@      "@     `h@      B@      @              4@     �K@       @      @      (@       @     �h@       @     @T@      "@       @       @      (@     �G@      @      @      J@      @     @X@      �?     �\@      ;@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @S�ƟH@�	           ��@       	                    �?���ŉ�@�            �@                           @�u�,�@J           (�@                            �?�7A!y�@           @{@������������������������       �F�,�h@�            `i@������������������������       �8�3әL@�             m@                            �?A`�Ɏ�@4           @������������������������       �@󙖎�?Y             b@������������������������       �|5$���@�            v@
                          �4@ȎAm
�@�           l�@                            �?d~9�_w@           �@������������������������       ��G`���@�            �p@������������������������       �AlO�r@^           ؁@                           @a��to<	@�           `�@������������������������       ��k�)��	@t           ؁@������������������������       �h�W�P@@(           �}@                           @i͂i)�@�           $�@                           �?'6���@           ��@                          �8@�F���@�           ��@������������������������       �x�8!�@&           �{@������������������������       �O�:d�E
@�             k@                           �?)=�$@^            `d@������������������������       ���T`3��?             <@������������������������       �~�V�g@O            �`@                          �7@��=�be@�            0q@                           @��2� @v             h@������������������������       ��Xt���?             G@������������������������       �ޡ$ˣ� @W            @b@                          �9@k�ak�@5            �T@������������������������       ���B���@            �E@������������������������       �Ѭ���@             D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     `t@     P�@      5@      M@     �{@     �X@     ��@     �j@     ��@     �u@      <@      $@     `m@     px@      @      C@      r@     �Q@     8�@     �c@      �@     @n@      4@      �?     �Q@     @_@      �?      @     �R@      .@     �u@      ;@     �k@      G@       @      �?      L@      K@               @     �F@      @     @\@      6@     �Z@      ?@      �?      �?      6@      @@              �?      3@       @     �J@      @     �N@       @                      A@      6@              �?      :@       @      N@      2@      G@      7@      �?              .@     �Q@      �?      �?      >@      &@     �l@      @      ]@      .@      �?                      (@      �?              (@      @     �S@              =@      @                      .@     �M@              �?      2@      @      c@      @     �U@      &@      �?      "@     �d@     �p@      @     �A@     �j@      L@     �z@     �`@     Pv@     �h@      2@             �N@      [@       @      @     @S@      &@     �p@     �H@     �f@     �R@                      3@      6@                      ?@      @      W@      5@     �G@      =@                      E@     �U@       @      @      G@       @     �e@      <@     �`@     �F@              "@     �Y@     �c@      @      =@      a@     �F@     �d@     �T@     �e@     �^@      2@      @      M@     �U@      @      1@     �T@      B@     �K@      P@      R@     �R@      0@      @     �F@      R@      �?      (@     �J@      "@     �[@      3@     �Y@     �G@       @      @     �V@     `d@      ,@      4@     @c@      ;@     �n@     �K@      j@     �Y@       @      @     @T@     `b@      &@      1@     �`@      8@      _@      J@     �`@      V@      @      @     �R@     @[@      $@      1@     �[@      4@     �U@     �A@     �[@     @R@      @       @      F@     @Q@      @      @     �T@       @     @Q@      ,@     @U@      K@      @      @      ?@      D@      @      $@      <@      (@      1@      5@      :@      3@       @              @      C@      �?              5@      @      C@      1@      7@      .@                      �?                              @              &@              &@      �?                      @      C@      �?              1@      @      ;@      1@      (@      ,@                      $@      0@      @      @      6@      @     �^@      @     �R@      .@       @               @      (@       @              "@      @      W@      �?      L@      @       @               @      @                                      9@              "@      �?       @              @      @       @              "@      @     �P@      �?     �G@      @                       @      @      �?      @      *@              ?@       @      3@       @                       @      @                      "@              2@              @      @                              �?      �?      @      @              *@       @      (@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ.�KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?$F,0�h@�	           ��@       	                    �?JE��vt@           h�@                          �<@e�� �>@�           x�@                           �?���خ@y           ��@������������������������       ����'sk@�            �k@������������������������       �_£�"D@�            0x@                          �=@Q9�e�
@             H@������������������������       �0e ���?             5@������������������������       �=mMm��@             ;@
                           �?�"��*Y@p           X�@                           �?�G��@�            pp@������������������������       �
�dd��@<            �Y@������������������������       ��Y/d@b             d@                           @D���ʳ@�            @t@������������������������       �����l�?�             m@������������������������       ��}��GC@<            �V@                          �5@�K��aU@�           ޤ@                           @��a�f�@r           `�@                           @8�x�Hg@�           ��@������������������������       ���K�I@_             d@������������������������       �w�=�P@q           ��@                           @]�]�S@�           Ѓ@������������������������       �es4;��@x           ��@������������������������       �@�ɟ&@*             O@                           �?�)X]=	@9           \�@                           @q/^!!
@�           x�@������������������������       �f�bw�	@h           ��@������������������������       ����f@6            �V@                           @?Y��aN@�           @�@������������������������       ����p��@�            �q@������������������������       �ֲ@�!@�            �v@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     ��@      ;@      Q@     |@     �T@     p�@      m@     p�@     pv@      :@             @W@     �d@       @      &@     �U@      @     �{@      D@     0r@     �Y@      @              E@     @V@      �?      "@     �F@      @      p@      ;@     @`@      H@                      E@     @U@      �?      @     �E@      @     @o@      7@      ^@     �@@                      <@     �@@      �?       @      0@      @      M@      0@     �E@      4@                      ,@      J@              @      ;@       @      h@      @     @S@      *@                              @              @       @      �?       @      @      $@      .@                              @                                      @              @      "@                                              @       @      �?      @      @      @      @                     �I@     �R@      �?       @      E@      �?     �f@      *@      d@     �K@      @              C@     �C@               @      ?@             �I@       @      M@     �A@      �?              *@      .@                      "@              :@      @      :@      "@      �?              9@      8@               @      6@              9@      @      @@      :@                      *@      B@      �?              &@      �?     ``@      @     �Y@      4@      @              $@      :@                       @      �?     @[@             �Q@      "@                      @      $@      �?              @              6@      @     �@@      &@      @      3@     `i@      y@      9@     �L@     �v@     �R@     ��@      h@     X�@      p@      6@      &@     �N@     `h@      "@      9@     @d@      <@     Pv@     �R@     `t@      \@      @      &@     �C@      \@      @      3@      ^@      .@      `@      P@     ``@     �U@      @       @       @      ,@              @      B@       @      ;@      (@      ?@      .@      @      @      ?@     �X@      @      .@      U@      *@     @Y@      J@      Y@     �Q@       @              6@     �T@      @      @      E@      *@     �l@      &@     `h@      :@       @              0@     �S@      @      @     �D@      &@      j@      $@      f@      2@                      @      @                      �?       @      4@      �?      2@       @       @       @     �a@     �i@      0@      @@      i@     �G@      f@     �]@     �h@      b@      .@      @     �T@     @[@      ,@      7@      W@     �A@     �I@     �Q@     �P@     �V@      *@      @     �Q@      Y@      *@      7@     �T@      =@     �F@     �E@      P@     @T@      "@       @      (@      "@      �?              "@      @      @      <@      @      $@      @      �?      N@     �X@       @      "@      [@      (@     �_@     �G@     @`@     �J@       @      �?      0@      D@       @      @     �G@      @     �R@      2@      J@      :@                      F@      M@               @     �N@      "@      J@      =@     �S@      ;@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ4��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @d,�4k@�	           ��@       	                   �5@�wK�%@�           ԥ@                          �1@�L�~�@�           ��@                           @�T�&��@#           }@������������������������       �b�:N[�@m            �e@������������������������       ���I���?�             r@                            �?�8iB�@�           l�@������������������������       ���g��p@           �z@������������������������       ��yC</Q@�           ��@
                           �?ܝ��n		@�           ��@                          �8@�W.)%@�            w@������������������������       �x�u��6@n            @h@������������������������       ��!QP�@o            �e@                          �<@!~�	@           h�@������������������������       ��k�wf	@�           p�@������������������������       �_��9��@\            �c@                           @�4���@�           |�@                           �?h.qGg�@           H�@                           �?�<�38	@�            �t@������������������������       �Բ�0�%@J            �^@������������������������       ��SA��%	@�            �i@                           �?�TW5@D            �@������������������������       ������@�            y@������������������������       �+���@E            �[@                           @�x�L�Y@�            `q@                          �1@�T���� @_            @d@������������������������       ��d|�?             ?@������������������������       �\���¡ @L            ``@                           @'�%z�@K             ]@������������������������       �w� ��?!             J@������������������������       ��Zv΅@*             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     Ps@     Ȁ@      :@     �I@     �z@     �U@     �@     �n@     ��@     �u@     �C@      &@     `l@      x@      0@     �@@      q@     �M@     h�@      e@     ��@     `n@      @@       @     �Z@     �l@      @      &@     @`@      1@     0�@     �P@     `w@     �\@       @       @      8@     �K@              @      >@      �?     @i@      0@     �Z@      :@               @      .@      8@                      ,@      �?      K@      .@      A@      0@                      "@      ?@              @      0@             �b@      �?      R@      $@                     �T@     �e@      @       @      Y@      0@     �s@     �I@     �p@     @V@       @              4@     �N@                     �G@      �?     �_@      4@     @]@      <@      @              O@     @\@      @       @     �J@      .@     �g@      ?@     �b@     �N@      @      "@     @^@     �c@      *@      6@      b@      E@     �l@     @Y@     �k@      `@      8@      �?      ?@     �I@       @       @      <@       @     @Z@      &@     �W@      =@      @              8@      <@       @      �?      .@             @P@      @     �G@      @       @      �?      @      7@              �?      *@       @      D@       @     �G@      6@      @       @     �V@     �Z@      &@      4@      ]@      A@     �_@     �V@      `@     �X@      1@      @     @R@     @X@      "@      2@     �U@      5@     �]@     �Q@      \@     �N@      *@       @      1@      "@       @       @      >@      *@      @      3@      0@      C@      @      "@     �T@     �b@      $@      2@     �c@      <@     �n@     �S@     �l@     �Z@      @      "@     �R@     �_@       @      .@      `@      ;@     �`@     �R@     `b@      W@      @      @     �B@     �I@      @       @      J@      .@      F@      1@      N@      ?@      �?              &@      "@      �?      @      4@      �?      9@       @      >@      &@              @      :@      E@      @      �?      @@      ,@      3@      "@      >@      4@      �?      @      C@     �R@      �?      @     @S@      (@      V@      M@     �U@     �N@      @      @     �@@     �K@      �?      @     �P@      (@     �M@      D@     �R@      G@      @              @      4@              �?      &@              =@      2@      (@      .@                      @      9@       @      @      <@      �?     @\@      @     @T@      ,@      �?              @      ,@                      4@      �?     @P@      �?     �J@       @      �?               @      @                                      0@              @                              @      @                      4@      �?     �H@      �?     �G@       @      �?               @      &@       @      @       @              H@       @      <@      (@                              �?              @      @              >@       @      &@      �?                       @      $@       @              @              2@              1@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��(JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @ǁ7�l@�	           ��@       	                   �8@@.	ڋ�@o           \�@                           �?N�٨�*@�           ��@                           @��@�           đ@������������������������       ���w�@           X�@������������������������       �d�Za�@�            `r@                          �1@J�r�f@%           �|@������������������������       �T^�g]k@7            @V@������������������������       �/�{�d�@�            Pw@
                           �?��� l�	@�           x�@                           �?^����	@0           �}@������������������������       �Sތ7	@g             c@������������������������       ����_�	@�            `t@                           @����V=@Y             b@������������������������       �������@=            �Y@������������������������       ���
���@            �E@                            �?�(�D@)           l�@                           @�`�ai@�            Py@                           �?����@�            �v@������������������������       ����]R$ @S            �^@������������������������       �����M�@�            @n@                           �?]�.�@             D@������������������������       �+O���?             .@������������������������       ��I��Xb�?             9@                           �?���yI*@+           �@                          �4@�)I<=@           �{@������������������������       �!�uk�?�             q@������������������������       �\-�}Ί@j            `e@                          �7@/؉fz9@           H�@������������������������       ���� @�           ��@������������������������       ��T�gı@�            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     (�@      A@     �M@     p}@     @U@     Ў@      l@     H�@     �u@      @@      1@     �j@     0t@      9@      F@      t@     �P@     �v@     �g@     px@     �m@      <@      &@     @d@      m@      0@      >@     @l@      <@     �s@     �]@     �s@     `a@      (@      &@     `a@     `d@      (@      :@     �d@      7@     �g@      T@     @k@     @X@      &@      @     @V@     @X@      &@      1@     ``@      .@     `d@     �H@     `g@     @Q@      "@      @      I@     �P@      �?      "@      B@       @      ;@      ?@      ?@      <@       @              7@     @Q@      @      @     �M@      @     �^@      C@     �W@      E@      �?              @      *@                                     �D@      "@      .@      @                      3@      L@      @      @     �M@      @     @T@      =@      T@     �A@      �?      @      J@     �V@      "@      ,@      X@      C@     �J@     �Q@     �S@      Y@      0@      @     �@@     �P@      "@      (@      S@      =@      A@      K@      K@     �V@      .@      @      &@      5@      �?      �?      <@      @      7@      *@      3@      7@      @      @      6@     �F@       @      &@      H@      9@      &@     �D@     �A@     �P@      $@              3@      9@               @      4@      "@      3@      0@      8@      $@      �?              @      6@               @      ,@       @      ,@       @      4@      "@      �?              .@      @                      @      �?      @       @      @      �?                      U@     @l@      "@      .@     �b@      3@     h�@      B@      z@     �[@      @              :@     �E@      �?       @      @@       @     @e@      $@     @T@      C@                      9@     �D@      �?              @@       @     @c@      @      S@      =@                              .@      �?               @      �?     @P@       @      8@      @                      9@      :@                      8@      �?     @V@      @      J@      6@                      �?       @               @                      0@      @      @      "@                                               @                      @      @      �?                              �?       @                                      "@              @      "@                      M@     �f@       @      *@     @]@      1@     0|@      :@     u@      R@      @              1@      R@              �?      4@       @     �i@      "@     @Y@      1@                      (@     �B@              �?      @             �c@      @     �I@      @                      @     �A@                      .@       @      H@      @      I@      $@                     �D@     �[@       @      (@     @X@      .@     �n@      1@     �m@     �K@      @              <@     �V@      @      @     �N@      .@     @j@      @     �e@      =@       @              *@      5@      @      @      B@             �A@      $@     �N@      :@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ,g+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?[9�v@�	           ��@       	                   �8@P��r	@�           ��@                            �?R�(ʙ@�           ��@                           �?���J:`@W           ؀@������������������������       �|Ge���@r            �e@������������������������       �3��-	@�            �v@                           �?����\�@K           X�@������������������������       �p�#�)�@~            �f@������������������������       �a|mfP�@�            `u@
                           �?�����V
@G           ��@                          �<@��&���@Y            �a@������������������������       �e��ߺ@5            �S@������������������������       ���$�@$             O@                           @:%At|
@�            Px@������������������������       �����	@4            @V@������������������������       �~��	��	@�            �r@                           �?"�w=,�@�           "�@                           �?7����@�            �@                          �<@b�"m_�@           �z@������������������������       ��N�_�� @�            �y@������������������������       �rD��*@             ,@                           @&6@�           �@������������������������       ��e�o�l@�            �o@������������������������       �Miߴ��@           �y@                           �?�W��@           $�@                            �?��Sʱ@�            �u@������������������������       ��Bk�=@v            @f@������������������������       �9�4@e            �e@                          �9@��ɇ|@&           X�@������������������������       ���E4�@�           (�@������������������������       �I�M��@m            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@      q@     ��@      >@     �Q@     �|@     �W@     P�@     �m@     ��@     pu@      >@      .@     `d@     �o@      2@     �G@     �o@     �L@      h@     �`@     �n@     �g@      8@      @      ^@      f@      &@      =@     �e@      ?@     �b@     �P@     �f@      ]@      @      @     @S@     �V@      @      "@     �T@      6@     �P@      @@     �X@     �H@      �?              7@      ?@               @      >@              A@      @      C@      "@              @      K@      N@      @      @     �J@      6@     �@@      9@     �N@      D@      �?      @     �E@     �U@      @      4@     @V@      "@     �T@     �A@     @T@     �P@      @      @      0@      <@      @      @     �A@      @      ?@      *@      3@      7@      �?              ;@      M@              0@      K@      @     �I@      6@      O@      F@       @      "@     �E@     �S@      @      2@     @T@      :@      F@      Q@      P@      R@      4@              .@      9@              $@      6@      �?      *@      (@      <@      ,@      �?              &@      *@              @      3@      �?       @      @      .@      @      �?              @      (@              @      @              @       @      *@      $@              "@      <@     �J@      @       @     �M@      9@      ?@      L@      B@      M@      3@      @      @      $@              @      "@      @      �?      *@      *@      &@      ,@      @      6@     �E@      @      @      I@      3@      >@     �E@      7@     �G@      @             �[@     @s@      (@      7@     @j@     �B@     H�@      Z@     �@     `c@      @             �K@     @a@      @      &@     �^@       @     0x@      H@     �n@     �R@      @              ,@     �E@              �?     �A@      @      k@      (@     �S@      8@                      $@     �E@              �?     �A@      �?     �j@      (@     @S@      5@                      @                                       @      @               @      @                     �D@     �W@      @      $@      V@      @     `e@      B@     �d@      I@      @              8@     �A@      �?       @      B@      @      H@      8@      L@      6@      @              1@      N@      @       @      J@      �?     �^@      (@     �[@      <@                      L@     @e@       @      (@     �U@      =@     `x@      L@     �t@     @T@      @              $@     �C@      �?              .@      @      c@      "@     �Y@      ,@       @              @      ?@      �?              @       @      Q@      @     �L@       @                      @       @                      (@      @      U@      @      G@      @       @              G@     ``@      @      (@      R@      8@     �m@     �G@     �l@     �P@      �?              9@     �]@      @      @      H@      3@     �k@      7@     �h@      G@      �?              5@      *@      @      @      8@      @      0@      8@      @@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�:0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�tqRBY@u	           ��@       	                    �?������@D           ��@                           �?�蒀�'@�           x�@                            �?��RSs�@"            }@������������������������       ����6�@�            �l@������������������������       �X�v��"@�            `m@                            �?�6�@d            �c@������������������������       ��V��@            �F@������������������������       ���@E             \@
                           @$�DK�{	@�           0�@                          �4@�%6AV	@F           �@������������������������       ��[a�� @L           ؀@������������������������       �R��Q��	@�           0�@                           �?.z񫯞	@x            `i@������������������������       ����T	@              N@������������������������       �κhX@X            �a@                          �2@iC�~�`@1           8�@                           @�v��@\           p�@                           �?���b���?�            �r@������������������������       ����$���?�             m@������������������������       �n�E��G @%            �P@                           @�3f�P�@�            0p@������������������������       �V �P�L@             i@������������������������       ��s�M@'             M@                           @����<@�           ��@                           @�ؑt4S@�           X�@������������������������       ��i4�K@�           ��@������������������������       ��#p���@
             3@                          �?@(����@�            Py@������������������������       ��B��@�            px@������������������������       ����v�t@	             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     `s@     @�@      B@     �I@     �y@     �U@      �@     `k@     0�@     �v@      ;@      2@      l@      t@      =@     �A@     �p@      O@     �x@     @f@     w@     �n@      8@       @      Q@     �R@      �?      @     �N@      @     �e@      :@     �a@     �L@      @       @      J@     @Q@      �?      @     �I@       @     �[@      6@     �Y@      F@      @       @      2@      @@              @      9@              H@      &@     �M@      =@      @              A@     �B@      �?      @      :@       @      O@      &@      F@      .@                      0@      @              �?      $@      @     @P@      @     �C@      *@                      @      @              �?       @       @      ,@              .@      @                      (@       @                       @      �?     �I@      @      8@      $@              0@     �c@     �n@      <@      <@      j@     �L@     �k@      c@     `l@     �g@      4@      ,@      a@     �k@      8@      :@     �e@     �H@      h@     @]@      j@     @e@      *@      @      ?@      T@      (@      @     @R@      @      `@     �E@      V@      N@      @      $@     @Z@     �a@      (@      3@     @Y@      E@      P@     �R@      ^@     �[@       @       @      5@      8@      @       @      A@       @      ;@     �A@      3@      4@      @      �?      @      @      @              "@      @       @      "@      @      *@       @      �?      ,@      4@               @      9@      @      9@      :@      ,@      @      @      �?     @U@     �p@      @      0@     �a@      9@     Ȃ@     �D@     P{@     �]@      @              *@      U@      �?      @      7@       @     �p@      @     �]@      B@       @              @      C@              �?      (@       @     �d@      @      L@      $@       @              @      9@              �?       @             �`@      @     �F@      "@       @               @      *@                      @       @     �@@              &@      �?                      @      G@      �?      @      &@             @X@       @     �O@      :@                      @     �B@                       @             @T@       @      I@      3@                      @      "@      �?      @      @              0@              *@      @              �?      R@     �f@      @      "@      ^@      7@     u@      A@     �s@     �T@      �?      �?     �F@      \@              @     �R@      *@     �n@      1@     �j@      K@      �?      �?      F@      \@              @      R@      "@      n@      *@     �j@      J@      �?              �?                               @      @      @      @      �?       @                      ;@      Q@      @      @      G@      $@     �V@      1@     @Z@      =@                      8@      Q@      @      @      G@      @     �V@      0@     �Y@      9@                      @                                      @              �?       @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>��<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�u��C@�	           ��@       	                   �2@�B���@b           "�@                           �?���'@!           `}@                          �1@6\^D�L@c            `c@������������������������       �>"�	��?7            @U@������������������������       �發"@,            �Q@                          �1@�;)�@�            �s@������������������������       �!�1� @i            �e@������������������������       ����l�@U            �a@
                           �?y���P�@A           �@                           �?R
vL8f@(           P}@������������������������       �r�Q��`@�            �u@������������������������       ��&�I�@M            �^@                           @gΟ��x	@           ��@������������������������       ����hl	@�           ܐ@������������������������       �����@g            �e@                            �?� ���@            ��@                          �4@E���@�            �x@                           @�<&��?~            �i@������������������������       �&����?v            @h@������������������������       �;z�0��@             $@                           �?N�}l+�@p            `h@������������������������       �J�.�@            �F@������������������������       �n�1�@V            �b@                          �6@ʤ����@2           ��@                           @���ּ2@@           ��@������������������������       �f�d�%�@{            `i@������������������������       ��a[-Bt@�           8�@                           @�1,�,0@�            py@������������������������       ���a��{@�            �q@������������������������       �Ч�$�@H             ^@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     pr@     H�@      @@     �K@      }@     �T@     0�@     `j@     @�@     0u@      9@      1@     �i@     `u@      7@      B@      t@      M@     Pw@     �d@     y@     �l@      3@       @      ?@     �N@      �?      @      Q@      �?     �^@      7@      [@     �F@      @              "@      2@              �?      &@      �?     �L@      �?     �H@       @                      @      ,@                      @             �D@              3@      �?                      @      @              �?      @      �?      0@      �?      >@      @               @      6@     �E@      �?       @     �L@             @P@      6@     �M@     �B@      @      �?      "@      8@      �?      �?      3@             �B@      ,@     �F@      7@              �?      *@      3@              �?      C@              <@       @      ,@      ,@      @      .@      f@     �q@      6@     �@@     �o@     �L@     `o@      b@     Pr@      g@      ,@      �?     �H@      W@      @       @     �E@      @     @Z@      4@     �Y@      F@      @      �?     �D@     �S@      @              =@       @      P@      1@     @R@     �B@       @               @      ,@               @      ,@       @     �D@      @      >@      @      �?      ,@     �_@     �g@      3@      ?@      j@     �J@     @b@      _@     �g@     �a@      &@      $@     �[@     �c@      3@      ?@     �f@     �F@      _@     �U@      f@     �_@      "@      @      0@      >@                      :@       @      6@      C@      ,@      .@       @      �?      V@     0q@      "@      3@      b@      9@     ��@      F@     pw@     @[@      @              ;@      D@               @      @@      @     �f@      &@     �Q@      >@                      @      .@               @      $@              _@      @     �@@      (@                      @      ,@                      $@             @^@      �?     �@@      $@                              �?               @                      @       @               @                      6@      9@                      6@      @     �L@       @      C@      2@                              "@                      @      @      5@      �?      @      @                      6@      0@                      2@       @      B@      @     �A@      ,@              �?     �N@     `m@      "@      1@      \@      4@     �{@     �@@      s@     �S@      @              <@     �d@      @       @      O@      (@     �v@      (@     @j@     �D@      @              &@     �D@                      *@      $@      R@      @     �B@      (@      @              1@      _@      @       @     �H@       @     @r@       @     �e@      =@      @      �?     �@@     �Q@      @      "@      I@       @      T@      5@     �W@      C@              �?      $@      I@      �?      "@      =@       @     �O@      *@      S@      ;@                      7@      4@       @              5@              1@       @      2@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���\�H@�	           ��@       	                    �?Z��ۯ�@�           <�@                           �?9|�5�Q	@           X�@                           �?7�0Lt@�           ��@������������������������       ��h*��@t            `e@������������������������       �A��JI@%           �|@                          �7@��×�	@~            �@������������������������       ����`��@|           p�@������������������������       ���ہ.
@            y@
                           �?�y�\2�@{           @�@                          �9@�֝�l�@p            �f@������������������������       �_�[M�8@^            �b@������������������������       ��^9�@             @@                          �3@
��ê�@           0y@������������������������       �j��@c            �a@������������������������       ����P@�            Pp@                          �4@`����@D           ��@                           @����^@N           ��@                          �2@�SN��@�            `j@������������������������       ��j��=��?Q            @^@������������������������       ��U;��@:            �V@                            �?�G��@�           (�@������������������������       �J��"��?`            �b@������������������������       �l팖��@c           x�@                           �?'����@�           ��@                          �5@r��N�]@�             y@������������������������       ��9�w}�@4             T@������������������������       ���'/� @�             t@                           @�c�?�#@           x@������������������������       �&��2�@�             u@������������������������       ��&��@"            �G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �t@     (�@      8@     �D@     p{@      U@     \�@     `l@     ��@     �u@     �D@      6@     @n@     Pr@      ,@      >@     `s@     �O@     �x@     �g@     �v@     �n@     �A@      6@      h@     `k@      *@      8@     `l@     �K@      m@     �a@     �p@     @h@      @@       @     �H@     �X@      �?      "@      W@      "@     @a@     �C@     @]@      Q@       @              .@      ;@                      (@              L@      @     �E@      &@       @       @      A@     �Q@      �?      "@      T@      "@     �T@      A@     �R@     �L@      @      4@      b@     @^@      (@      .@     �`@      G@     �W@     �Y@      c@     �_@      8@      *@     �V@     @T@      @      @     �P@      (@     @S@      I@     �Z@     @R@      &@      @      K@      D@      "@       @     @Q@      A@      1@     �J@     �F@     �J@      *@             �H@     �R@      �?      @     �T@       @     `d@      H@     �X@     �I@      @              2@      *@                      1@              S@      @      D@      &@      �?              ,@      @                      *@             @R@      @      >@      &@                      @       @                      @              @       @      $@              �?              ?@     �N@      �?      @     �P@       @     �U@     �E@      M@      D@       @              @      8@               @      &@             �G@      1@      ;@      "@                      :@     �B@      �?      @     �K@       @      D@      :@      ?@      ?@       @             �V@      l@      $@      &@      `@      5@     `�@     �B@     Pz@     �Z@      @             �F@     �Z@      @      �?     �H@       @     @{@      2@     `k@     �C@                      6@      ;@                      @       @      X@      @     �G@      @                       @      *@                                      Q@      @      8@      @                      ,@      ,@                      @       @      <@       @      7@      �?                      7@      T@      @      �?     �E@             @u@      *@     �e@     �@@                      @      0@                      $@             �U@              <@      @                      4@      P@      @      �?     �@@             �o@      *@      b@      ;@                     �F@     @]@      @      $@      T@      3@      k@      3@     @i@     �P@      @              ?@      P@              @      C@      $@     �\@      @     �Y@      :@      @               @      0@                      "@      @      8@              1@       @      @              =@      H@              @      =@      @     �V@      @     �U@      8@      �?              ,@     �J@      @      @      E@      "@     @Y@      .@     �X@     �D@       @              @     �H@       @      @      A@       @      W@      &@     @X@     �B@                      "@      @      @               @      �?      "@      @       @      @       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJI�GhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����-@�	           ��@       	                    �?�1}�U�@           h�@                          �;@�n *�@8           `}@                          �5@��R�@           Py@������������������������       ��3�P�@�            `o@������������������������       �g��`@l            @c@                           �?zmF�@(            @P@������������������������       ��UQ�@             7@������������������������       ��ȷ^�X@             E@
                          �2@YMc�l	@�           �@                            �?�,朙i@~             i@������������������������       �	--�7�@!             K@������������������������       �y�F@]            `b@                           @:o�	@K           ؍@������������������������       ��38>|@�            �l@������������������������       ��c�6��	@�           ��@                          �4@fS�C�@�           ޡ@                          �1@:��x@�           �@                            �?���-@           �y@������������������������       �	L�
3% @E            �Y@������������������������       ��Ρa:@�            @s@                          �3@��h�@�           8�@������������������������       �#���@W           ��@������������������������       ���RQ�(@�            �n@                          �7@��"��@�           ��@                           @��e-@;           �@������������������������       �Udv�@�            s@������������������������       ��8�_�t@x             i@                           @p�zBf@n           ��@������������������������       �x9�#��@�            �u@������������������������       �$[���@�            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �t@     �@      7@     �K@     @{@      S@     �@     �j@     ��@     �w@      6@      2@     `g@     `k@      .@      @@     �n@      D@     `o@     �_@     �p@      j@      3@      �?     �F@     �T@      �?      $@     �J@      @     �[@      9@     �W@     �D@      �?             �A@      S@      �?      @     �G@      @     @[@      4@     �T@      :@      �?              ,@      F@              @      5@      @     �T@      &@     �K@      1@                      5@      @@      �?      �?      :@              :@      "@      <@      "@      �?      �?      $@      @              @      @      �?       @      @      (@      .@              �?      @      @                      @              �?              @      @                      @      @              @      �?      �?      �?      @      @      (@              1@     �a@      a@      ,@      6@     �g@      B@     �a@     �Y@     @e@      e@      2@      @      8@      ;@      �?      �?      D@              C@      "@      ;@      ;@       @              @      @                      *@              0@      �?       @      @              @      2@      4@      �?      �?      ;@              6@       @      3@      8@       @      (@     �]@     @[@      *@      5@     �b@      B@     �Y@     @W@     �a@     �a@      0@      @     �D@      4@      @      �?     �F@       @      $@      4@      D@      A@      @       @     @S@     @V@      "@      4@     �Z@      <@      W@     @R@     �Y@     �Z@      (@             @b@      t@       @      7@      h@      B@     8�@      V@     H�@     �e@      @              H@     �d@      @      &@     �R@      @     0@      C@      r@     @T@                      @     �M@              @      2@             �h@      ,@     �U@      9@                              1@              �?      @             �K@      @      &@      $@                      @      E@              @      ,@             �a@      $@     �R@      .@                      E@      [@      @      @     �L@      @     �r@      8@     @i@      L@                      >@     �R@       @      @      C@      @     �j@      $@      c@     �A@                      (@      A@       @      @      3@      @     �U@      ,@      I@      5@                     �X@     `c@      @      (@     @]@      >@     @q@      I@      m@      W@      @              F@     @V@       @      �?     �I@      3@     �b@      @     �\@      ?@      �?              4@     �C@       @      �?     �A@      ,@     @Z@      @     �P@      2@                      8@      I@                      0@      @     �E@              H@      *@      �?              K@     �P@       @      &@     �P@      &@      `@      G@     �]@     �N@       @              G@     �C@              "@     �D@      $@     �R@      <@      P@      B@       @               @      ;@       @       @      9@      �?     �J@      2@      K@      9@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?=ep(2@�	           ��@       	                   �;@=�>,�+	@�           D�@                           �?r�X�@%           L�@                            @f�ʨp@�             w@������������������������       ���2�+@�            @k@������������������������       ������@`            �b@                           �?����)	@6           �@������������������������       �oW���@�            �u@������������������������       � ǳ�y	@\            �@
                           �?TB8��	@�            �o@                            �?�H���@5            @Q@������������������������       �tAZ��@             3@������������������������       ��h�UJ�@&             I@                          �>@�u��	@z             g@������������������������       �W!����	@O             ^@������������������������       ���Z'1@+            @P@                          �5@���t�@�           p�@                           @�iO@�           ��@                          �1@���\4�@X           t�@������������������������       �S��J @           �z@������������������������       ��o��ٷ@T           ��@                           �?C\���1@8            @X@������������������������       ��kr�Ε@            �C@������������������������       �m<U�u@$             M@                           @*=w�@#           Ћ@                           @��/�[@�           ��@������������������������       �śZDԤ@f           p�@������������������������       �P�p�)1@~            �h@                           �?����Y�@?            �Y@������������������������       �<�@             A@������������������������       �F��YxE@)             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     ��@      A@     �D@     P{@     �S@     ��@      h@     p�@     �w@     �@@      0@     �e@      p@      6@      9@     @m@      H@     �i@     @[@      n@     �h@      9@      "@     �a@      k@      *@      1@     �i@      A@      g@     @W@     �k@     @a@      8@              B@     @P@      �?      @     �B@      �?      V@      2@     @T@      ?@      @              6@      ?@               @      ;@      �?      G@      @     �M@      2@      @              ,@      A@      �?       @      $@              E@      (@      6@      *@              "@     �Z@      c@      (@      *@     @e@     �@@     @X@     �R@     `a@     �Z@      2@              8@     �S@      @      "@     @P@      @      J@      2@      I@      F@      @      "@     �T@     �R@      "@      @     @Z@      =@     �F@     �L@     @V@     �O@      ,@      @      >@     �C@      "@       @      ;@      ,@      6@      0@      4@     �N@      �?      �?      @      &@              �?       @       @      (@      @       @      3@                              @                      @              @       @      @      �?              �?      @      @              �?      @       @       @      �?      @      2@              @      :@      <@      "@      @      3@      (@      $@      *@      (@      E@      �?      @      4@      (@      @      @      *@      $@      "@      @      @      :@               @      @      0@      @      �?      @       @      �?      @      @      0@      �?       @     @_@     `u@      (@      0@     `i@      ?@     h�@      U@     ��@     �f@       @             �G@     `l@      @      &@     @V@      0@     ��@     �C@     @w@     @T@      @             �E@     �j@      @      @     �U@      ,@     ��@      A@     0v@     �P@      @              1@      J@              @      (@             `j@      @     �[@      (@       @              :@     `d@      @      @     �R@      ,@     �t@      ;@     �n@      K@      �?              @      (@              @       @       @      @@      @      1@      .@      @              @                      @       @       @      &@      �?      @       @       @              �?      (@                                      5@      @      (@      @      �?       @     �S@     �\@      @      @     �\@      .@     �i@     �F@     @i@     @Y@       @       @      K@      Z@      @      @     �X@      *@      h@      ?@     @g@     @X@       @       @      F@      Q@              @     �S@      @     @d@      2@     �a@      P@       @              $@      B@      @      �?      3@      @      >@      *@     �F@     �@@                      8@      &@      �?              0@       @      ,@      ,@      0@      @                      &@       @                      @              @      @      @                              *@      "@      �?              "@       @      @      $@      *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�w�ChG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����8?@�	           ��@       	                    �?�$�-2	@           ��@                          �<@\R�d@<           �~@                          �3@5�q�R�@            {@������������������������       �Q�+���@q            �e@������������������������       �jÊ�ɛ@�            p@                           �?t<��7@(             M@������������������������       ���x�@             1@������������������������       �t&KY��@            �D@
                          �1@� �	�	@�           �@                            �?�?�;@G            @]@������������������������       �ⴿ{j@)            @Q@������������������������       �܊&�N&@             H@                           �?�E��	@�           �@������������������������       �O�B��h	@�             u@������������������������       ����z=�	@�           ��@                           �?� '���@�           ̡@                          �2@�pO��@�           X�@                            �?���C�?�            @r@������������������������       ����	�5 @[             a@������������������������       ��j>���?^            `c@                           @�����x@            p|@������������������������       �Ĩ��r@�            �t@������������������������       ���/�h�@Q            �^@                          �1@lDF	@�           �@                           @�O�@2@�             o@������������������������       ���1�K@(             O@������������������������       �~�=���?z            @g@                           @]1��J�@7           �@������������������������       �sz@,-+@�           ��@������������������������       �����@w            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     @r@     P�@      ?@     �I@     P~@      Q@     ��@     �k@     ��@     �v@      8@      8@     �d@     �l@      8@      @@     `p@     �B@     �n@      a@      p@     �i@      4@      �?      K@      Q@      �?      @     �M@      @     @\@      :@     @Y@      I@      @      �?     �G@      N@      �?      @     �I@      @      [@      7@      X@      @@      @              &@      6@                      8@      @      H@       @      D@      .@              �?      B@      C@      �?      @      ;@              N@      .@      L@      1@      @              @       @              @       @              @      @      @      2@                      @      @                      �?              @              �?       @                       @      @              @      @              �?      @      @      0@              7@     �[@      d@      7@      9@     `i@      >@     ``@     �[@     `c@     �c@      1@      �?      "@      0@      �?              *@      �?      =@      @      ;@      ,@              �?       @      0@                      @      �?      &@      @      ,@      "@                      �?              �?              @              2@      @      *@      @              6@     �Y@      b@      6@      9@     �g@      =@     �Y@     @Z@      `@     �a@      1@      "@      ;@     @R@      *@      @     @P@      @      ;@      A@      8@     �E@      "@      *@     �R@     �Q@      "@      3@     @_@      7@     �R@     �Q@      Z@     �X@       @             �_@     `t@      @      3@     �k@      ?@      �@     �U@     ��@     @c@      @              ;@     �Z@                      K@      @     pt@      (@      g@      >@      �?              $@      5@                      2@              d@      @      P@      *@      �?               @      ,@                       @             �Q@              ;@      "@                       @      @                      $@             �V@      @     �B@      @      �?              1@     @U@                      B@      @     �d@       @     @^@      1@                      .@     �M@                      8@      @     �`@      @     �S@      *@                       @      :@                      (@              A@      @      E@      @                      Y@     �k@      @      3@      e@      :@     �y@     �R@     �w@      _@      @              @     �A@               @       @             �Z@      $@     �Q@      (@                       @      1@                      @              0@      @      $@      @                       @      2@               @      @             �V@      @     �N@      @                      X@      g@      @      1@      d@      :@     �r@      P@     Ps@      \@      @             �Q@     �d@      @      1@      a@      5@     �p@      F@     �p@      W@      �?              :@      4@      @              9@      @     �B@      4@      C@      4@       @�t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�h�UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@M�ʱ�6@�	           ��@       	                    @��푟]@�           ��@                           �?zE$�_B@E           �@                          �0@�[tiLU@�            �r@������������������������       �"UD>@            �A@������������������������       ����p�a@�            �p@                          �3@��1���@�           ��@������������������������       ���2�]@#           �|@������������������������       �yB�(�@a             a@
                           @�H�]Z@D           (�@                          �2@¨��9@�            �@������������������������       ��
?4.�?            {@������������������������       �z
�(4a@�            �n@                           �?$j#���@�            p@������������������������       �$}4�@X            �a@������������������������       �k��?ma@D             ]@                           �?��U@!           F�@                           �?2��qg@	@u           @�@                           �?N���)O@�            �p@������������������������       �]5�Yu@K            �]@������������������������       �R�ij�
@Z             c@                           �?����	@�           І@������������������������       �E�Y�B�@�            �n@������������������������       ����	@8           `~@                          �6@%�a��k@�           �@                           �?�BE_@�            �v@������������������������       ��j�Ƭ�@}            @h@������������������������       ����ՍA@v             e@                          �;@xYփ�@�           ��@������������������������       ���{�w@C           ��@������������������������       ���Mq��@v            @f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �q@     h�@      >@     �M@     P~@      S@     p�@      i@     ȉ@     �w@      9@       @     �W@     �m@      $@      .@     �h@      2@     (�@      T@     Px@     �d@      @       @     �M@     �\@       @      (@     �b@      "@     �i@      N@     `d@      \@      @              <@     �C@               @     �C@      �?     �V@      $@      N@      =@      �?              �?      @                      (@              ,@       @       @      �?                      ;@      B@               @      ;@      �?      S@       @      M@      <@      �?       @      ?@     �R@       @      $@     �[@       @     �\@      I@     �Y@     �T@      @       @      9@      N@      @      "@     @R@      @      Y@     �C@      S@     �Q@      �?              @      .@      @      �?     �B@      @      ,@      &@      ;@      *@      @              B@     �^@       @      @     �H@      "@     �y@      4@     @l@     �K@       @              6@      Y@              �?      <@      @     Ps@      *@     �d@      ?@                      ,@     �P@                      ,@      �?      k@       @      Z@      ,@                       @     �@@              �?      ,@      @     @W@      &@     �O@      1@                      ,@      6@       @       @      5@      @      Y@      @     �M@      8@       @              @      ,@       @       @      &@      @     �K@      @      ?@      (@                      "@       @                      $@             �F@       @      <@      (@       @      *@     �g@     t@      4@      F@     �q@      M@     �v@      ^@     @{@     �j@      2@      (@     �_@      d@      (@     �A@     �c@      :@     �T@      R@     �e@     @`@      ,@       @      G@     �F@              (@      @@              ;@      *@      L@      B@      �?       @      7@      1@              &@      (@              @      "@      9@      ,@                      7@      <@              �?      4@              6@      @      ?@      6@      �?      $@      T@      ]@      (@      7@     @_@      :@      L@     �M@      ]@     �W@      *@      @      ,@      F@      @       @      E@      @      :@      ,@      H@     �@@      @      @     �P@      R@      @      .@     �T@      6@      >@     �F@      Q@     �N@      $@      �?     @P@      d@       @      "@     @`@      @@     `q@      H@     �p@      U@      @              *@     �L@               @     �J@      &@     @]@      "@     �U@      ,@      �?              @      7@               @      C@      "@      P@      @      C@      "@                      @      A@                      .@       @     �J@      @      H@      @      �?      �?      J@     �Y@       @      @     @S@      5@      d@     �C@     @f@     �Q@      @      �?     �@@      R@      @      �?      I@      .@      a@     �A@     @a@      J@      �?              3@      ?@      �?      @      ;@      @      8@      @      D@      2@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ 0i4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@>	��ц@�	           ��@       	                    �?v�����@g           �@                           @0�7}�@�            �@                            @�1b^U@�            �t@������������������������       �k�%���@�            �i@������������������������       �����@S            �_@                           @��=V2�?           �y@������������������������       �`���T @=            �Y@������������������������       ��x��\�?�            0s@
                           @�9-�+@�           0�@                          �1@u�ȋ�@�           ��@������������������������       ��O�,�@x            `g@������������������������       �U����	@h           Ё@                          �1@7��b�@�           ��@������������������������       ��QI���?x             f@������������������������       �(ض�i@4           `~@                          �<@���@S           d�@                           �?.`7��V@�           `�@                           �?�4�΢@�            @y@������������������������       �~sF�1q@z             j@������������������������       �0�@��@x            `h@                          �7@���^�@�           �@������������������������       ���69@           �x@������������������������       �P�/��	@�           ��@                           @�uQI�@�            t@                           @z����@�            �p@������������������������       ���2	�@�            �n@������������������������       ���[�@             9@                           @L{�w�@!             I@������������������������       �(�l&>�@             7@������������������������       ��8I���@             ;@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     @t@     �@      <@      O@     0{@     @U@     `�@     �l@     ��@      w@      ?@      *@     �]@     �r@      &@      ?@      i@      <@     ��@      Y@      ~@     �e@      (@             �D@     @X@      @      �?     �H@      @     pt@      1@      d@     �C@      @              :@     �B@      @      �?     �A@              U@      ,@     @X@      ?@      @              &@      5@      @              8@              G@       @     �Q@      3@      @              .@      0@              �?      &@              C@      @      ;@      (@                      .@      N@                      ,@      @     `n@      @     �O@       @                      @      4@                      @      @     �H@              4@      �?                      $@      D@                      $@             @h@      @     �E@      @              *@     @S@     `i@       @      >@      c@      9@     �v@     �T@      t@      a@      "@      *@      J@     �[@      @      7@     @Z@      .@     �`@     �R@     �^@     �W@      @      �?      (@      C@                      1@             �H@      4@      ?@      3@              (@      D@     @R@      @      7@      V@      .@     �U@      K@      W@     �R@      @              9@      W@      �?      @     �G@      $@     �l@      "@     �h@      E@      @              @      0@              @       @             �T@              K@       @                      6@      S@      �?       @     �C@      $@     @b@      "@     �a@      A@      @      @     �i@     q@      1@      ?@     @m@     �L@     �q@     @`@     s@      h@      3@      @     @d@     �k@      $@      5@     �g@      D@     @p@      Y@     q@      `@      3@              F@      N@      @      �?      G@      @     �V@      .@     @[@      :@      @              6@      ;@      @      �?      <@             �M@      @      G@      0@                      6@     �@@                      2@      @      @@       @     �O@      $@      @      @     �]@      d@      @      4@      b@     �A@      e@     @U@     �d@     �Y@      .@      �?     �M@     �S@              "@     �H@      *@     �P@      3@      L@     �C@       @      @     �M@     �T@      @      &@      X@      6@     �Y@     �P@      [@      P@      @      �?      F@      J@      @      $@     �E@      1@      5@      >@      @@      P@              �?     �E@     �D@      @       @     �@@      0@      $@      >@      :@     �L@              �?     �B@      D@      @       @      :@      0@      $@      >@      6@      I@                      @      �?                      @                              @      @                      �?      &@      �?       @      $@      �?      &@              @      @                      �?      @               @      @              @              �?                                      @      �?              @      �?      @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Ԙ`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?v��F@�	           ��@       	                    �?������@"           ��@                           @���+j�@�           ��@                            �?�x���@�            �s@������������������������       �	c�>�@n             d@������������������������       �z��o� @]            �c@                          �5@�J�h9- @�            �u@������������������������       ��cF@_��?�             n@������������������������       ���}@<            �Y@
                            �?[xLe8@�           ��@                           �?��y<-@�            �t@������������������������       ��
t���@b             c@������������������������       �j�5�@o             f@                           @�ҽ@�            �p@������������������������       ��,u@c            `b@������������������������       �v�4���?P            �]@                          �1@B����@�           ��@                           @y��۠@�            pv@                           �?7�D�E@#            �O@������������������������       ��S�8��?	             .@������������������������       ���Z�P@             H@                            �?���x@�            �r@������������������������       ����Vއ@n             f@������������������������       ������@P             ^@                          �:@y_���p@�           �@                           @K�i^�,@�           �@������������������������       ���_�9	@�           ��@������������������������       ��O aD@           ؈@                           @���ʽ@           `{@������������������������       �s���h�@           @z@������������������������       �u���#�?             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�         @     �t@     H�@      =@      K@     �|@     @S@     ��@     @k@      �@     �w@      @@             @V@      e@      @      *@     �[@      (@     �|@      D@     Pq@     �S@      @             �B@     �S@      @      (@      L@       @     q@      .@     �a@      B@      �?              ;@      C@      @       @     �C@      @     �W@      (@     @P@      9@      �?              "@      6@       @      @      .@      �?     �H@       @      @@      .@      �?              2@      0@      �?      �?      8@      @     �F@      @     �@@      $@                      $@     �D@              @      1@      �?     `f@      @     �S@      &@                      @      =@              @      @             �a@      �?      H@      @                      @      (@                      (@      �?      C@       @      >@      @                      J@     �V@      �?      �?      K@      @      g@      9@     �`@      E@      @              9@      P@      �?      �?      9@       @      V@      $@     �T@      9@      @              .@      ;@              �?      3@             �@@      @     �A@      .@      �?              $@     �B@      �?              @       @     �K@      @      H@      $@      @              ;@      :@                      =@       @     @X@      .@     �I@      1@       @              7@      3@                      8@       @      ?@      $@      6@      0@                      @      @                      @             �P@      @      =@      �?       @       @     �n@      x@      9@     �D@     �u@     @P@     0�@     @f@     �~@     �r@      9@       @      7@      I@              @      :@             �_@      1@      S@     �A@                      ,@       @                      �?              5@      @      $@      "@                                                                       @      @      �?      @                      ,@       @                      �?              *@      @      "@      @               @      "@      H@              @      9@             @Z@      &@     �P@      :@               @       @      ;@               @      (@              P@      @     �C@      7@                      @      5@               @      *@             �D@      @      ;@      @              @     �k@     �t@      9@     �B@      t@     @P@     �z@      d@     �y@     pp@      9@       @     �d@     @r@      4@      >@     `n@      J@      w@     �`@     v@     �f@      4@      �?     �[@      d@      .@      :@      f@     �C@      a@     �\@      c@      ]@      1@      �?     �J@     ``@      @      @     �P@      *@      m@      2@      i@     �P@      @      @      M@      E@      @      @     @S@      *@      L@      =@      O@      T@      @      @      I@      E@      @      @     �Q@      *@      L@      ;@      O@      T@      @      �?       @                              @                       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�8�/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @X4q�m@�	           ��@       	                    �?ML���@x           ��@                          �;@Ǚ'uY�@�           �@                           �?¼#�ֿ@s           8�@������������������������       �Nq#�Bd@           `z@������������������������       �嚆e�@e             d@                            �?����H@7            �V@������������������������       ��=�@             9@������������������������       �����a@*            @P@
                          �9@6����l	@�           Ę@                          �1@�F�q��@�           ��@������������������������       ��<OG�@b             d@������������������������       ��Q�	@v           �@                           �?)v���
@�            �x@������������������������       ���>�9w	@c            �c@������������������������       ���m��	@�             n@                           �?{�a[r�@           ܙ@                            �?��a��� @f           P�@                           @X��|� @O            �^@������������������������       �X�Җ��?$            �M@������������������������       �`����?+             P@                          �2@�v	�� @           �z@������������������������       �t�b~�?o            �f@������������������������       �3���_@�            @o@                          �7@Y۬�'�@�           4�@                          �1@�#�}/�@
           ؉@������������������������       �C��� @z            �i@������������������������       ��R)�g@�           h�@                           @M�#�@�             q@������������������������       ���4m�@             G@������������������������       �
�\?B@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     `�@      D@      I@     `~@     @T@     x�@     �i@     Ј@     `w@      @@      1@     �l@     �t@     �@@     �@@     �u@     �P@     @u@      e@     �x@     �p@      ;@             @Q@      Z@       @      "@     �U@       @     �c@      8@     �b@     �N@      @             �K@     @V@       @      @      Q@      @      c@      5@     @a@      H@       @              F@     �R@       @      @      I@       @     �Y@      4@     �T@      C@       @              &@      ,@                      2@       @      I@      �?     �K@      $@                      ,@      .@              @      3@      @      @      @      $@      *@      @               @      "@                       @      @                       @      @      @              (@      @              @      1@              @      @       @      $@              1@      d@     �l@      ?@      8@     Pp@     �M@      g@      b@     �n@      j@      6@       @     �\@      g@      9@      2@      k@     �@@     �b@     �Z@     �h@     �_@      &@              &@      8@      �?              2@              D@      1@      @@      1@               @     �Y@      d@      8@      2@     �h@     �@@     �[@     @V@     �d@     @[@      &@      "@      G@      G@      @      @      F@      :@      A@     �C@     �G@     �T@      &@      @      3@      7@      @       @      4@      $@      @      $@      (@     �C@      @      @      ;@      7@       @      @      8@      0@      ;@      =@     �A@     �E@      @      �?     �Q@     �k@      @      1@     @a@      ,@     ؃@      C@      y@     @Z@      @              7@     @P@      �?             �A@       @     `q@       @     �]@      7@      �?                      *@      �?              &@      �?      O@      �?      9@      "@                               @                      �?              @@              "@      "@                              @      �?              $@      �?      >@      �?      0@                              7@      J@                      8@      �?      k@      @     @W@      ,@      �?              "@      *@                      @             @\@      �?     �A@      @      �?              ,@     �C@                      3@      �?     �Y@      @      M@      $@              �?      H@     �c@      @      1@     �Y@      (@     Pv@      >@     �q@     �T@      @              A@      _@      @      "@      N@      &@     pr@      *@     �l@      F@       @               @      >@               @      (@             �T@      @     @Q@      @                      @@     �W@      @      @      H@      &@     �j@      "@      d@     �C@       @      �?      ,@     �@@      �?       @     �E@      �?      O@      1@      K@      C@       @      �?       @       @      �?      @      @              "@      �?      @      @                      (@      9@               @     �B@      �?     �J@      0@      H@      @@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�99FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @z���`@�	           ��@       	                   �4@�aE_�@�           p�@                           �?j��J@A           x�@                           �?]�(�6�@}           h�@������������������������       �7�.s�;@�            �j@������������������������       ��?�2;�@�            �w@                           @���/h@�             t@������������������������       �Lk�@:o@�            �m@������������������������       �$�s��@/             U@
                          �9@1�D��|	@@           ��@                           �?�ғ0	@�           H�@������������������������       ��`�%�<	@�           �@������������������������       �����@r             e@                           �?�#l+��	@F            �@������������������������       �f��w��	@
           �y@������������������������       ��ju�m�@<            �X@                           @�w6�@#           D�@                           �?Vf
8`'@�           4�@                            �?�
c�%B @�            @w@������������������������       �6r;ˠ	�?9            �V@������������������������       ��} Yk @�            �q@                          �6@�����/@�           Ȉ@������������������������       ��q���@d           �@������������������������       �����\r@�             k@                          �4@��c��@K            �@                           @S�Ct@�             n@������������������������       �r��L�@�            @l@������������������������       ��[� -��?             ,@                           @j��O�@�            @q@������������������������       �MzZ�v�@�            �o@������������������������       ���I�@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     �@      @@      L@     @@      X@     ��@      l@     Ȉ@     �s@      9@      5@      k@     �t@      >@     �C@     �u@     @R@     �w@     @g@     �w@     @j@      1@      @     �N@     �a@      @      &@     �^@      0@     �k@     @P@     `f@      T@      @      @     �G@     @T@      @      @      V@      ,@     ``@      E@     �Z@      M@      @       @      ,@      B@      @      �?      B@      @      L@      2@      6@      3@              @     �@@     �F@      �?      @      J@      $@     �R@      8@     @U@     �C@      @              ,@      N@              @      A@       @     @V@      7@      R@      6@                      &@      A@              @      @@              P@      ,@      L@      5@                      @      :@                       @       @      9@      "@      0@      �?              ,@     `c@     �g@      9@      <@      l@     �L@     �c@     @^@     `i@     @`@      *@      @      Z@     �\@      0@      6@      b@      8@     �[@     �P@     �_@     �P@      "@      @     �U@     �V@      0@      2@      ^@      0@     �R@     �J@     @Z@      I@       @              2@      8@              @      9@       @     �B@      ,@      5@      0@      �?      "@     �I@     @S@      "@      @      T@     �@@      H@      K@     @S@      P@      @      "@      F@     �P@      "@      @      O@      9@     �A@      E@      L@      L@      @              @      $@              �?      2@       @      *@      (@      5@       @               @     @T@     �j@       @      1@      c@      7@     ��@     �C@     �y@     �Y@       @       @     �L@     �a@               @      Y@      (@      ~@      6@     pq@      M@      @              0@     �I@                      6@       @     �g@       @      S@      (@                              (@                       @              J@              *@      @                      0@     �C@                      ,@       @     `a@       @     �O@      @               @     �D@      W@               @     �S@      $@     r@      4@     `i@      G@      @              4@     �R@              @     �H@       @     `n@      @     �a@      ;@      @       @      5@      2@              @      =@       @      G@      *@      O@      3@      �?              8@     �Q@       @      "@     �J@      &@     �b@      1@     �`@      F@      @              &@      6@      �?      @      :@             �X@       @      K@      5@      �?              "@      5@      �?      @      9@             �X@       @     �I@      ,@      �?               @      �?                      �?                              @      @                      *@      H@      �?      @      ;@      &@     �I@      .@     �S@      7@      @              "@     �G@              @      5@      $@      I@      (@     �R@      7@                      @      �?      �?              @      �?      �?      @      @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ8K�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@:����J@�	           ��@       	                    @,/�N��@a           2�@                           �?��3@�           ��@                          �3@��kG@           �{@������������������������       �=���j@�            `r@������������������������       ������@`            �b@                           �?&�ʏ�@�           ��@������������������������       ��pn@*            ~@������������������������       ����%��@�             j@
                           @ӡ�l@�@�           ��@                            �?B:�%�:@�            0q@������������������������       �h�Gご�?'            �O@������������������������       ��޴�@w            �j@                            �?p��"�@           ��@������������������������       �4蘕5��?f            �b@������������������������       �%$i/@�           �@                           �?M���]�@?           ��@                           �?3|-��@)           `}@                          �<@R�W[�@�            �n@������������������������       �����k@r            @g@������������������������       ���Ԅ�@#             M@                          �>@�{'�@�            @l@������������������������       �ќK��Z@�            `j@������������������������       �/p3O�@
             .@                           @e�� i	@           h�@                           �?���V��	@            �@������������������������       ��nd��@+            �O@������������������������       �ROs�]	@�           �@                            �?��
	7@	           �y@������������������������       ��<h�(@I             \@������������������������       ���T�f@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     `r@     �@     �@@      I@     �}@     �R@     �@      i@     ��@     �v@     �A@       @     �W@     @s@      3@      =@     �l@      ?@     ��@     �S@     �}@     �f@      1@       @     �N@     @d@      2@      7@     �d@      5@     `o@      P@     �j@     �`@      ,@      @      3@      Q@      "@      @     �S@      &@     �W@      A@     �O@     �K@      �?      @      *@     �D@       @              H@      @     �Q@      7@      E@      F@      �?              @      ;@      @      @      >@      @      8@      &@      5@      &@              @      E@     �W@      "@      1@     �U@      $@     �c@      >@      c@     �S@      *@      @      C@      M@      @      "@     �Q@      "@      W@      4@     �X@     @P@      *@              @      B@       @       @      1@      �?      P@      $@      K@      *@                      A@     @b@      �?      @     @P@      $@     �}@      .@     �p@      I@      @              @      H@                      *@      "@     @]@      @      P@      *@      @              �?      *@                                      @@       @      &@      @                      @     �A@                      *@      "@     @U@      �?     �J@      "@      @              =@     �X@      �?      @      J@      �?     0v@      (@      i@     �B@                      @       @              �?      $@             �W@      �?      6@      "@                      9@     �V@      �?      @      E@      �?     @p@      &@     @f@      <@              1@     �h@      m@      ,@      5@     �n@     �E@     �r@     @^@      t@     �f@      2@      �?      F@      R@      @      @      M@       @     @]@      2@      ]@      ?@      @      �?      D@     �E@              @      A@      �?     �@@      *@      K@      3@       @      �?     �@@      <@               @      7@      �?      ?@      $@     �G@       @       @              @      .@               @      &@               @      @      @      &@                      @      =@      @              8@      �?      U@      @      O@      (@      �?              @      =@      @              2@             �T@      @     �M@      "@      �?              �?                              @      �?      �?              @      @              0@     `c@      d@      $@      1@     �g@     �D@     �f@     �Y@     �i@     �b@      .@      .@     �]@     @\@      @      ,@     ``@      C@     �Q@      U@     �[@     �]@      ,@      @      "@      $@              @      *@                      @      $@      @      �?      &@     @[@     �Y@      @       @     �]@      C@     �Q@     �S@      Y@     �\@      *@      �?     �B@      H@      @      @     �L@      @     �[@      3@     �W@     �@@      �?              1@      (@                      $@             �@@      �?      7@      0@              �?      4@      B@      @      @     �G@      @     @S@      2@     �Q@      1@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�q�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@.���3#@�	           ��@       	                    �?;Ƶ
@l           x�@                          �1@0��|"@e           @�@                           �?͕"����?�            `o@������������������������       �cT�L�� @,             Q@������������������������       ��||��?s            �f@                          �4@o��ߊ?@�           h�@������������������������       ����&�(@�            `w@������������������������       ��Z�@�            pu@
                          �4@��kg%@           П@                           @f/��I@�           `�@������������������������       �WU���@�           ��@������������������������       �J)�6@n           (�@                           @М�� �@           ��@������������������������       �ö}#��@;           �@������������������������       �5�@�             v@                          �<@���b�G	@N           h�@                           �?�ӱ�]�@�           ��@                           @�\���*
@�            Ps@������������������������       ��b%b	@�            �h@������������������������       �PX�ݞ�	@E             \@                           �?��q�W�@�            �q@������������������������       ���JF"��?*            �Q@������������������������       ���74��@�             k@                           @Ci��W<	@�            �s@                           �?a@U'	@�            �l@������������������������       ��s�^��@*            @Q@������������������������       ��;�f�@o             d@                           @��<*�@4            �T@������������������������       �^�>���@            �C@������������������������       �0ɞ�+W@             F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �p@     ��@      <@     �Q@     �z@      Q@     ȏ@     @k@     �@     Pw@      >@      @     �g@     �{@      0@     �J@     �s@      D@     Ћ@     @^@     ��@     �o@      .@             �F@      `@      @      @      P@      @      y@      =@     �l@      M@      �?               @      >@                      *@             @b@      @      I@      @      �?                      (@                      @              ?@      @      *@       @                       @      2@                      @             �\@      �?     �B@       @      �?             �E@     �X@      @      @     �I@      @     �o@      8@     @f@      K@                      3@      G@               @      1@      �?     �a@      0@     @Y@      @@                      8@      J@      @      @      A@      @     �\@       @     @S@      6@              @     �a@     �s@      (@     �G@      o@     �A@     �~@      W@     0{@     �h@      ,@       @     @Q@     �d@      @      3@      `@       @     �t@      M@     `p@      _@       @       @     �E@     �U@      @      *@      W@      @      ^@      I@     @^@     �T@       @              :@     �S@      �?      @      B@      @      j@       @     �a@      E@               @     �R@     `c@      @      <@      ^@      ;@     @d@      A@     �e@     @R@      @       @      L@     �Z@      @      ;@      T@      .@     �O@      ;@      R@      J@      �?              2@      H@              �?      D@      (@     �X@      @     @Y@      5@      @      $@      T@     �]@      (@      1@     �\@      <@     �_@     @X@     �e@     �]@      .@      "@      E@     �S@      @       @     �O@      "@     �Z@      Q@     �`@      N@      *@      "@      ?@      E@      @      @     �H@      @     �A@      D@     �E@      =@      *@      @      ;@      <@      @      @      B@       @      3@      5@     �@@      &@      @       @      @      ,@      @      �?      *@      @      0@      3@      $@      2@      @              &@      B@              @      ,@       @     �Q@      <@     �V@      ?@                              $@                              �?      7@       @      =@      @                      &@      :@              @      ,@      �?      H@      :@      O@      9@              �?      C@     �D@      @      "@     �I@      3@      5@      =@      C@      M@       @      �?      <@     �@@      @       @      ?@      1@      &@      ;@      4@     �H@       @               @      $@              @      $@              @      @      &@      .@       @      �?      4@      7@      @      @      5@      1@       @      5@      "@      A@                      $@       @      @      �?      4@       @      $@       @      2@      "@                              @      @      �?      @       @       @       @      @      @                      $@      �?                      .@               @              (@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$OphG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @N�7��o@�	           ��@       	                   �2@�����@�           ��@                           �?K��@=           �}@                           �?���=��@�             r@������������������������       �5��W@]            �`@������������������������       �m9���@o             c@                           �?��Ŋy�@q            `g@������������������������       �b�D���?&            �O@������������������������       �mZk��(@K             _@
                          �;@<Y�/n	@c           �@                           �?��gY	@�           �@������������������������       ����x�F@            �y@������������������������       �#[� m	@�           ��@                           �?T�t�\
@�             t@������������������������       �^�Lo�#	@B            �[@������������������������       ��ҥ��	@�             j@                           �?=t�@1           ��@                          �4@���Z� @n           ��@                          �1@��ӱo��?�            0v@������������������������       ���k�?f            @c@������������������������       ���|��?y             i@                           @&2�+�@�             j@������������������������       �5�U��@:             S@������������������������       �Ziyfޜ@U            �`@                           @�&"}H�@�           �@                           @k��@�            �@������������������������       �m$]9� @^            �b@������������������������       �Sx���@�           ��@                          �4@�.&\�G@�            Ps@������������������������       ����Z@W            �_@������������������������       �sH~@v            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     �r@     ȁ@      ?@      J@     �}@      O@     �@     @k@     H�@     �y@     �A@      ;@     @m@     pu@      7@      E@      u@      J@     �w@     �f@     Pu@     pq@      @@      �?      9@     @P@       @      �?      P@       @     @a@     �D@     �T@      J@       @      �?      5@      C@       @      �?      I@      �?      P@      5@      I@     �B@       @      �?      @      *@                      2@              E@      ,@      <@      &@      �?              ,@      9@       @      �?      @@      �?      6@      @      6@      :@      �?              @      ;@                      ,@      �?     �R@      4@      @@      .@                      �?      @                       @              >@              2@      @                      @      6@                      (@      �?      F@      4@      ,@       @              :@      j@     `q@      5@     �D@      q@      I@      n@     �a@     0p@     `l@      >@      (@     �e@     `m@      1@      >@      m@     �B@     `k@     @]@     �k@     �c@      5@             �N@     �L@      @       @      G@             �[@      7@     �R@      >@      @      (@     @\@     @f@      *@      <@     `g@     �B@      [@     �W@     `b@     �_@      1@      ,@     �A@     �E@      @      &@     �C@      *@      5@      8@     �B@     �Q@      "@       @      (@      3@              @      0@              @      @      (@      5@      @      @      7@      8@      @      @      7@      *@      0@      3@      9@     �H@       @              O@     @l@       @      $@     @a@      $@     8�@      B@     @y@     �`@      @              &@     �T@      �?              ?@      @     �p@      @      a@      8@                      @     �@@                      2@              h@      @     @V@      ,@                       @      2@                      (@             @W@              :@      @                      @      .@                      @              Y@      @     �O@      &@                      @     �H@      �?              *@      @     @R@       @      H@      $@                      @      .@                      @      @      >@      �?      (@      @                       @      A@      �?              $@             �E@      �?      B@      @                     �I@      b@      @      $@     �Z@      @     �u@      ?@     �p@      [@      @             �C@      [@      �?      @      Q@      �?     �q@      2@      g@      L@       @              .@      8@              @      0@              I@      @      9@       @                      8@      U@      �?      �?      J@      �?     �m@      ,@      d@      H@       @              (@      B@      @      @     �C@      @      O@      *@     �T@      J@      �?              @      0@      @       @       @              C@       @      C@      *@                      @      4@       @      �?      ?@      @      8@      &@      F@     �C@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJZ��ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?P#<W5@�	           ��@       	                    �?l����*@           �@                          �8@Pe��-@�           ��@                          �7@;c��x)@L           H�@������������������������       ���"48�@-           �}@������������������������       ��n�\�@             G@                            @�r`�@I            �\@������������������������       �^�$@)             Q@������������������������       ���kFq�@             �G@
                          �6@B���}�@m           P�@                          �2@f�E�9@�            �x@������������������������       �E4Ib@~            `i@������������������������       ��P��z@z            �h@                           �?�z��@u            `g@������������������������       �i�@C             [@������������������������       ��뙋�R@2            �S@                           @c�gܼ/@�           �@                           �?4h��	@�           ��@                           �? u�K7�@M             `@������������������������       ��Y|cT�@             C@������������������������       �m\<+\6@9            �V@                           �?,�ˀbI	@o           ��@������������������������       �Xy����	@�           ��@������������������������       �������@�            �w@                           @f�d2�@�           l�@                          �<@#g�␸@�           �@������������������������       ��"�nf@�           �@������������������������       ��{9n@&             Q@������������������������       �G����@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        *@     pr@     �@     �@@     �H@     �z@     �V@     ��@      g@     ��@     �w@      C@             @S@      f@      @       @      \@      $@     0z@      >@     �s@     �P@      @              ?@     �X@       @       @     �J@      @      n@      4@     `a@      B@      �?              7@     �R@       @      @     �G@      @      k@      $@     @]@      5@      �?              1@     @P@      �?      @      F@      @     `i@      $@      Z@      5@      �?              @      "@      �?      �?      @              *@              *@                               @      9@              @      @       @      8@      $@      6@      .@                      @      6@                               @      (@      @      (@      &@                      @      @              @      @              (@      @      $@      @                      G@     @S@       @             �M@      @     `f@      $@      f@      >@      @             �@@     �I@                     �@@             `a@      @     @_@      *@      �?              @      1@                      7@             �U@      @     �L@       @      �?              :@      A@                      $@              J@      �?      Q@      @                      *@      :@       @              :@      @      D@      @      J@      1@       @              $@      .@                      5@              *@      @      ?@      &@       @              @      &@       @              @      @      ;@      �?      5@      @              *@     @k@      w@      =@     �D@     �s@      T@     ȁ@     `c@     �@     �s@      A@      (@     �b@     �k@      6@      :@     �j@     @P@     �g@     �_@     �m@     �j@      ?@      @      (@      *@               @      A@      @       @      0@      *@      0@      @              �?       @                      @      @              @       @      $@      @      @      &@      @               @      =@       @       @      (@      &@      @               @     @a@      j@      6@      2@     �f@      N@     �g@     �[@      l@     �h@      :@       @      Z@     �a@      2@      2@      c@      H@     �\@     �T@      b@     �b@      :@              A@     �P@      @              =@      (@     �R@      ;@      T@      H@              �?      Q@     �b@      @      .@      Z@      .@     �w@      =@     Ps@     @Y@      @      �?      P@     �b@      @      .@     �Y@      &@     pw@      ;@     @s@      Y@      @      �?      K@      b@      @      .@      T@      &@     �v@      ;@     �r@      V@      @              $@      @      �?              6@              "@              "@      (@                      @              @               @      @      @       @      �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?C}�kP@�	           ��@       	                    @E�z<a�@           |�@                           �?��7�v�@�           �@                           �?�=��6@2           `}@������������������������       ����=@v            �f@������������������������       �d��@�            r@                          �<@����^�@|            �i@������������������������       �<C�k�@t             h@������������������������       ����aM@             *@
                           �?hܻ���@l           ��@                            @����C@�            �t@������������������������       � �fl��@�            pq@������������������������       ��Uu@���?#            �K@                            �?��ސy�@�            �m@������������������������       �e�L8�� @&            �M@������������������������       ��c�T��@t            `f@                           @����@�           Ԥ@                           �?���ic	@�           ��@                           �?��>8	@O            @a@������������������������       �~����t@7            �V@������������������������       ����N%�@             H@                          �3@8�N�F	@�           `�@������������������������       ��A�U@           �y@������������������������       �4����	@�           �@                          �6@w_�1�@�            �@                           @D�#	�I@�           X�@������������������������       �+'{�@�           ��@������������������������       ��g�L@	             *@                           @򰲫�r@�            �w@������������������������       ���)T� @�            �o@������������������������       ��.��o|@R             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     s@     (�@      =@     �K@     �{@      U@     ��@     �h@      �@     �w@      ;@      �?     @Z@     �e@      @      $@      X@      &@     {@      A@     �q@     @U@      @      �?     �U@     @Z@      @      "@     �N@      @     �e@      ;@     �a@     �K@      @      �?      L@     �U@      @      @      G@       @     @Z@      8@     �V@      F@      @      �?      ,@      >@                      2@              K@       @     �G@      *@       @              E@      L@      @      @      <@       @     �I@      6@      F@      ?@      @              ?@      3@              @      .@       @      Q@      @     �I@      &@      �?              ?@      2@              @      $@       @     �P@      @      H@      "@                              �?                      @              �?              @       @      �?              2@     �Q@       @      �?     �A@      @     @p@      @     �a@      >@                      (@      A@              �?      :@      @     @d@      @     @S@      ,@                      $@      ?@                      :@      @      `@      @      P@      &@                       @      @              �?                     �@@              *@      @                      @      B@       @              "@       @     �X@      @     @P@      0@                              @       @              @       @      ?@              (@      @                      @      ?@                      @             �P@      @     �J@      (@              5@      i@     `y@      7@     �F@     �u@     @R@     p�@     �d@      �@     @r@      4@      4@      a@     �o@      7@      @@     �m@     �N@     �l@      a@     �k@     @i@      2@      @      1@      0@              @      :@      @      @      1@      4@      4@      @      @      $@      "@                      1@      @      @      *@      1@      &@      @              @      @              @      "@      �?      @      @      @      "@              0@     �]@     �m@      7@      ;@     �j@     �L@     �k@      ^@     @i@     �f@      .@      @      5@      N@       @      �?     �K@      @     �Z@     �B@     @P@     �I@      @      (@     �X@      f@      5@      :@     �c@     �J@     �\@     �T@      a@     ``@      &@      �?      P@      c@              *@     �[@      (@     �t@      ;@     `r@     �V@       @              ?@      Y@              $@     �K@      @     @p@      @     �h@     �H@       @              ?@     �X@               @      J@      @     0p@      @      h@     �H@       @                       @               @      @       @      �?              @                      �?     �@@     �J@              @     �K@      @     �Q@      5@     �X@     �D@              �?      6@     �A@                     �D@      �?      L@      &@     @Q@      1@                      &@      2@              @      ,@      @      ,@      $@      =@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ	�_XhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�a��E@�	           ��@       	                   �<@��2洴@�           ��@                          �2@M�	$e@�           �@                           �?�S.[@.           �}@������������������������       ���b���@�            �t@������������������������       ��[�5{g@_            `b@                          �8@}u!��@�           ��@������������������������       ��*�K]@�           ��@������������������������       ���?�	@�            �w@
                           �?%��!	@�            �o@                          �?@m2om�W@0            �S@������������������������       �!Jb�@%             P@������������������������       ���i���@             ,@                           �?z*�X�W	@q            �e@������������������������       ����u�@)             N@������������������������       �,	�Z�	@H            �\@                            @��P��@1           �@                            �?����=@�           �@                          �7@	�Ϧ�@N           ��@������������������������       �%6D_j@�           �@������������������������       ��aɩs@v             f@                          �5@{x��%9@6           �|@������������������������       �Bn�y�@�             r@������������������������       ��zG���@t            �d@                          �3@m+7��@�            �p@                          �0@C2BC��?K            �[@������������������������       ���x�G��?
             .@������������������������       �n���0�?A            �W@                           @l�u	�@b            �c@������������������������       �&�2B��@[             b@������������������������       �X��*�@             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      s@     ��@      >@      P@     P}@      S@      �@     @i@     ��@     `w@      7@      3@     �m@     Ps@      7@      F@     �u@     �L@     @v@     �d@     Py@     �p@      2@      *@     �j@      q@      4@     �B@     s@      G@     �u@     �`@     �w@     �i@      .@      @     �B@     �P@              �?      S@      @     �_@      =@     @U@      G@       @      @      >@      G@              �?     �N@      @     �R@      2@      N@      =@       @              @      5@                      .@             �I@      &@      9@      1@               @      f@     �i@      4@      B@     �l@     �E@     �k@      Z@     �r@      d@      *@      @     �`@     `c@      .@      <@     �d@      9@     �d@     �O@     `n@     @_@      @      @     �D@      J@      @       @      P@      2@     �K@     �D@     �J@      B@      @      @      9@     �A@      @      @      D@      &@      $@      @@      8@     �L@      @              @       @               @      $@              @      1@       @      6@       @              @      @              �?      @              @      0@      @      6@       @               @      �?              �?      @              �?      �?      @                      @      4@      ;@      @      @      >@      &@      @      .@      0@     �A@      �?      @      @      0@      �?              *@      @              @      @       @              �?      0@      &@       @      @      1@      @      @      &@      *@      ;@      �?      �?      Q@     �k@      @      4@      _@      3@      �@     �B@     0z@     �[@      @      �?      N@      h@      @      .@     �Z@      3@     ��@     �B@     �t@     �W@       @              B@     @]@      @      "@     �N@      1@     Pv@      9@     �n@     �R@                      6@     �V@      @       @     �E@      (@     �t@      *@     �h@      G@                      ,@      :@              �?      2@      @      7@      (@     �H@      <@              �?      8@     �R@      @      @     �F@       @     @f@      (@     �U@      5@       @              *@     �F@              @      0@             �a@      @     �J@      &@       @      �?      &@      >@      @       @      =@       @     �B@      @      A@      $@                       @      <@              @      2@             @Z@             @U@      .@      @              @      ,@                      @              H@              C@       @                               @                                      &@              �?      �?                      @      (@                      @             �B@             �B@      �?                      @      ,@              @      .@             �L@             �G@      *@      @               @      &@              @      .@             �K@              F@      *@                      �?      @                                       @              @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�p(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?QKv�ia@�	           ��@       	                    �?`oL��@�           �@                           �?Yuo��@3           �~@                            @D,�@x             i@������������������������       �4���y@X            �a@������������������������       ���NriV @              M@                           �?�ېMV@�            0r@������������������������       �d}�Gl@W            @a@������������������������       ��XٱA~@d             c@
                           @��w��%@�           p�@                          �8@�0<$�@$           �|@������������������������       ���� � @�            `x@������������������������       ��4�~�@)            �P@                           �?u_!�o]@�            `p@������������������������       ��]�Gq@V            `a@������������������������       �e�j�O�@N            �^@                          �4@�c�=@�            �@                           @2�c8f�@�           \�@                            @���@�             n@������������������������       �o�侱�@d            �e@������������������������       �8%��;>@*            �P@                          �1@.���N�@P           8�@������������������������       �nT�p�O@�            �p@������������������������       ���b2�@�           Є@                           @$��D�	@�           �@                           @�K.���	@Y           P�@������������������������       �>���C	@           p{@������������������������       ��a���	@@           ��@                           @}��x@]           x�@������������������������       ����C0@�            �w@������������������������       �ioj�A0@q            @f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     @t@     ؀@      >@     �M@     �|@     @S@     ��@     `l@      �@     �v@      >@             @V@     @e@      @      "@     @[@      @     �z@     �C@     0p@     �U@      @              L@     �S@               @     @Q@      @     �Y@      7@     �W@     �J@      @              6@      :@                      ?@             �O@      @     �C@      $@       @              5@      0@                      ;@              C@      @      7@      "@       @              �?      $@                      @              9@      �?      0@      �?                      A@     �J@               @      C@      @      D@      0@     �K@     �E@      �?              2@      :@              @      0@      @      1@      (@      2@      4@      �?              0@      ;@              �?      6@              7@      @     �B@      7@                     �@@     �V@      @      �?      D@      @     �t@      0@     �d@      A@       @              <@      L@                      7@      @     �k@      &@     �W@      4@      �?              <@      H@                      5@      �?     @h@      @     @T@      *@                               @                       @       @      :@      @      *@      @      �?              @     �A@      @      �?      1@              [@      @     �Q@      ,@      �?              @      2@              �?      *@              Q@       @      9@      @                              1@      @              @              D@      @      G@      @      �?      0@     `m@     w@      9@      I@     �u@     �Q@     ��@     �g@     �@     q@      9@      @     �S@     �b@      (@      ,@     `a@      "@     t@     �P@     �p@      Z@      @      @      9@      9@      �?      @      >@      @     �G@      2@      M@      5@      @              3@      (@               @      :@       @      @@      ,@     �G@      0@      @      @      @      *@      �?      �?      @      �?      .@      @      &@      @                     �J@     @_@      &@      &@     @[@      @      q@      H@     `j@     �T@      @              *@      F@              @      8@              V@      @     @S@      *@                      D@     @T@      &@       @     @U@      @     @g@     �D@     �`@     �Q@      @      $@     �c@     `k@      *@      B@     �j@      O@     �m@     �^@      q@      e@      2@      $@      \@      d@      (@      >@      c@     �H@      Z@     �W@     �^@     �[@      *@      @     �C@     �J@      @      $@     �S@      >@      L@      B@      P@      O@       @      @     @R@      [@      "@      4@     �R@      3@      H@     �M@      M@      H@      &@             �F@      M@      �?      @      N@      *@     �`@      ;@     �b@     �M@      @              <@      C@              �?      C@      @     @[@      (@      [@      B@      @              1@      4@      �?      @      6@      @      :@      .@      E@      7@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ\��fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @x`��@�	           ��@       	                   �2@�%�=�@e           �@                            �?��FY<@/           �}@                           �?@���	@Z            �b@������������������������       ��ؒ.E�@7            @X@������������������������       �\N���@#             K@                           �?.��]0@�            0t@������������������������       ���d�@@T            �^@������������������������       �q5u7�I@�             i@
                            �?�O�egl	@6           ��@                           @���L	@4            ~@������������������������       �ù$��	@�            @r@������������������������       �U��Ee%@o            �g@                          �?@�w��S	@            �@������������������������       �s�-	@�           �@������������������������       �X@��}�@%            �P@                          �4@��8@�@=           �@                            �?vb�͵�@F           ��@                          �1@c�ĩI�?�            �i@������������������������       ���K3��?5            �R@������������������������       �����?Q             `@                           �?i��4�(@�           ��@������������������������       �4�+e�v @�            �q@������������������������       ��b��nU@            }@                           @~�V�m@�           H�@                          �7@p�	I��@�           H�@������������������������       ��9�P%f@�            �t@������������������������       ���#o��@�            �u@                          �5@i��)�@:             X@������������������������       ���7�g�?             .@������������������������       ���_�@2            @T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     `�@      @@     @Q@     @}@     �U@     8�@     @k@     `�@     �t@     �E@      ,@     `j@     `u@      4@     �J@     �t@     @P@     �u@     �e@     �v@     �l@      ?@       @      ?@     �R@      �?              Q@      @     ``@      ?@      V@     �D@      @              @      <@                      4@      @      H@      &@      ;@       @      �?              @      1@                      3@       @      9@      "@      1@      @      �?              �?      &@                      �?      �?      7@       @      $@      @               @      :@     �G@      �?              H@             �T@      4@     �N@     �@@       @       @      $@      1@      �?              ?@              ;@      @      ,@      ,@                      0@      >@                      1@              L@      ,@     �G@      3@       @      (@     �f@     �p@      3@     �J@     �p@      O@     �j@     �a@     0q@     �g@      <@      @      L@     �K@      �?      1@     @R@      &@      Q@      H@     �U@      H@      (@      @      @@      A@              "@      F@      &@     �F@      (@      M@     �@@       @              8@      5@      �?       @      =@              7@      B@      =@      .@      @      @      _@     �j@      2@      B@     �g@     �I@     `b@     @W@     �g@     �a@      0@      @     @Z@     �i@      ,@      ?@     �f@      H@     @b@     @V@     �f@     �`@      0@       @      3@      @      @      @      "@      @      �?      @      @      @                     �Y@     �n@      (@      0@      a@      6@     h�@      G@     z@     �Y@      (@             �K@     �]@      @      $@      H@      @     @z@      0@     �l@     �G@      @              @      3@              �?      @             @]@      @     �C@      0@                              @              �?       @              I@      �?      &@      @                      @      ,@                       @             �P@       @      <@      &@                      I@     �X@      @      "@      F@      @     �r@      *@      h@      ?@      @              0@     �A@               @      "@             �a@      @     @R@      @      @              A@      P@      @      @     �A@      @     `d@      $@     �]@      :@                     �G@      `@      @      @      V@      3@      i@      >@     @g@      L@      "@              A@     �]@      @      @     �T@      1@      f@      3@     @e@     �J@      �?              4@     @R@      @      �?      ?@      "@     @Y@      @     �S@      *@      �?              ,@      G@              @     �I@       @      S@      0@     �V@      D@                      *@      "@      @              @       @      8@      &@      0@      @       @                                                      �?      @              @      �?      @              *@      "@      @              @      �?      5@      &@      *@       @      �?�t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJluShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@[�V_�-@�	           ��@       	                   �1@ןe��@�           ��@                           �?+l|��@�           ��@                           @#<M,@�            �s@������������������������       �f�:��@�            �m@������������������������       ��T�8@,             S@                           @���.�(@�            �s@������������������������       ��{販�@i            �b@������������������������       �Q��R��?h             e@
                           @!Y3E�@�           ��@                           @�Z?b�E@�           (�@������������������������       ��\A�@t           �@������������������������       ��d��l�@i            `d@                           �?ŏz*ė@"           0}@������������������������       �%d.��?m             g@������������������������       ���o��@�            �q@                           @Bg���@"           4�@                           �?�?�[MN	@H           ��@                           �?xr6�	@�           ȏ@������������������������       ���|�@�            �t@������������������������       ��w�4��	@�           X�@                           �?e���@�            `t@������������������������       ��Qׄy@V            �`@������������������������       ��s��'.@p            �g@                            �?F�J ��@�           ؆@                          �5@q� 8h�@y            �g@������������������������       ��w+�]'�?            �A@������������������������       �FO@�V@d            @c@                          �7@��yJ?�@a           ��@������������������������       ����@�            0q@������������������������       �XA�@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �q@     ��@      =@     �J@     0z@     �S@     (�@     �m@     @�@     pv@      >@      @     �V@     �n@      @      1@     @e@      .@      �@     @U@     �z@     �`@      @      �?      8@     �T@      @      @     �G@      �?     �p@      5@     @b@      ?@              �?      "@      E@      @      @      9@      �?     �a@      (@     �M@      0@                      @     �A@      @              6@             �Z@      @     �H@       @              �?       @      @              @      @      �?     �A@      @      $@       @                      .@      D@              �?      6@              `@      "@     �U@      .@                      &@      :@              �?      1@             �D@      @      B@      &@                      @      ,@                      @              V@       @     �I@      @               @     �P@     �d@      @      (@     �^@      ,@      w@      P@     �q@     �Y@      @       @     �H@     @\@      @       @     @Y@      (@      c@     �K@     `d@      S@      @       @      ?@      U@      @      @      V@      &@      _@      A@     �_@     @P@      @              2@      =@               @      *@      �?      =@      5@     �B@      &@       @              1@     �I@      �?      @      6@       @      k@      "@     �]@      :@                       @      .@                      @             @Z@      @      F@      @                      "@      B@      �?      @      1@       @      \@      @     �R@      7@              $@     `h@     `t@      6@      B@      o@     �O@     Pv@      c@     �y@     @l@      8@      $@     �b@     `l@      2@      >@     @f@      F@     @c@     �^@     `l@     `d@      6@      $@     �^@     �e@      2@      7@     ``@      ?@      [@     @X@      c@     �`@      4@              >@     �J@      �?      @      G@      @      K@      7@     �Q@      D@      @      $@      W@      ^@      1@      1@     @U@      <@      K@     �R@     @T@      W@      *@              :@      K@              @     �G@      *@      G@      9@     �R@      ?@       @              "@      &@              @      8@      @      =@      (@      <@      *@      �?              1@     �E@              @      7@      "@      1@      *@     �G@      2@      �?             �G@     �X@      @      @     �Q@      3@     `i@      ?@     @g@     �O@       @              7@      7@      @              1@      @      M@      @      E@      *@                              @                      @              &@              0@       @                      7@      4@      @              ,@      @     �G@      @      :@      &@                      8@      S@      �?      @      K@      .@      b@      9@      b@      I@       @               @     �H@      �?      @      4@      &@      W@      @      Q@      .@      �?              0@      ;@              �?      A@      @     �J@      4@      S@     �A@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�9�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����V@�	           ��@       	                    �?�p]E�@M           ��@                           �?���=>	@�           ��@                           �?f�WA�V@3           @~@������������������������       ��]HG۶@u             f@������������������������       �2@�D�@�            0s@                          �:@���E��	@�           �@������������������������       ��M]�{	@           p�@������������������������       �@:�4�	@�            �n@
                           �?�P�i,#@b           P�@                            �?���1�J@^            �a@������������������������       ���\@             I@������������������������       �y�� ��@?             W@                           �?<�xU�@           �y@������������������������       ���ؙ��@g             c@������������������������       ��m1u��@�            @p@                          �5@BzT$6@s           �@                           �?f�<l�I@�           ��@                            �?�v"�@�           ��@������������������������       �^���}�@�             v@������������������������       ���j�S�@�            �n@                           @3�M@Q           ��@������������������������       �C�Q�t��?�            �w@������������������������       ����U��@\             c@                          �<@_fn��@�           x�@                            @8+�[g@\           8�@������������������������       ��:���@           �{@������������������������       ��Ġ�j� @=            �Z@                            �?�yMf @@             Z@������������������������       �"���+~@$             L@������������������������       ��+з@             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     @�@      B@      N@     �~@     �P@     0�@     �i@     X�@     �v@      @@      3@     �j@     @t@      <@     �D@     �t@     �I@     �v@     �d@     �t@     �l@      :@      3@     �f@     �m@      :@      B@     �p@      C@     `l@      ]@     @l@      f@      5@       @     �L@     �R@      @      @     @Q@      @     �Y@      <@     �U@     �H@       @       @      2@      ;@                      8@              H@      @     �A@      .@      �?             �C@     �G@      @      @     �F@      @     �K@      5@      J@      A@      �?      1@      _@     �d@      7@      >@      i@      A@      _@      V@     `a@      `@      3@      @     �W@     �`@      2@      :@      d@      9@     �Y@     �K@     �]@      V@      1@      $@      =@      @@      @      @     �C@      "@      5@     �@@      4@      D@       @              @@     �U@       @      @      P@      *@     �`@     �I@     �Z@      K@      @              @      3@              �?      $@             �I@      @      E@      @      @                      "@              �?      �?              .@              3@      �?      @              @      $@                      "@              B@      @      7@      @                      <@     �P@       @      @      K@      *@      U@      G@     @P@      H@      �?               @      ;@                      6@      @      ;@      *@      :@      8@      �?              4@      D@       @      @      @@      "@     �L@     �@@     �C@      8@               @     @U@     �l@       @      3@     �c@      0@     �@      D@     �y@      a@      @             �C@     �c@      @      @     �R@      @      @      &@     @p@     �Q@      @              8@     �Q@       @      @     �K@       @     �o@      @     �`@     �D@       @              $@      C@      �?      @     �B@      �?     �b@      @     �U@      4@       @              ,@     �@@      �?      @      2@      �?     �Z@             �G@      5@                      .@     �U@      �?      �?      3@      @     `n@      @     �_@      =@      @              @     @P@      �?      �?      @      @     `g@       @     �V@      1@                       @      5@                      *@      �?      L@       @     �B@      (@      @       @      G@     �Q@      @      (@     �T@      $@      f@      =@     @c@     �P@      �?       @      C@     �N@      @      $@      J@      $@     �c@      ;@     `a@      I@      �?       @      C@      K@      @      @      F@      $@      Z@      :@     �[@      G@      �?                      @       @      @       @              J@      �?      =@      @                       @      $@               @      ?@              4@       @      .@      0@                      @      @                      .@              @       @      (@      (@                      @      @               @      0@              .@              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�e{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�U}m�P@�	           ��@       	                   �1@V�L���@u           ��@                           �?�Po�,@�            �p@                           �?s�(Q�@?            @W@������������������������       ��_�lO�?             >@������������������������       ����d�V@*            �O@                          �0@�-g���@o             f@������������������������       �ƎY�]@            �I@������������������������       ��I-@Q            @_@
                            �?���f2	@�           ��@                          �<@�]#�G	@�           ��@������������������������       �,&ǈ��@<           x�@������������������������       �����@G             Y@                           �?'5i��@D           ؋@������������������������       ���e��	@�           ��@������������������������       ���/u^@�            `i@                           @��:/@:           8�@                          �2@2��v_@�           ��@                           @����l��?
           �y@������������������������       ���Ri��?�            �h@������������������������       ��t�i@�            �j@                           @�M��Y@�           P�@������������������������       ��^�y�@�           ��@������������������������       �y>�@             8@                           @�s���@W           @�@                           @d�A�A@@           @�@������������������������       ���p���@           �{@������������������������       ��.���;@3             S@                           �?�
�W��	@             @@������������������������       ��$��� @	             *@������������������������       �,l��ۛ@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     ȁ@      :@     �K@     �}@     �T@     �@     `j@     ؇@     �t@      =@      8@     �k@     `r@      ,@     �F@     Pt@     �Q@     �x@      e@     �u@     @m@      :@       @      3@      @@              @      5@      �?      Y@      0@      H@      ;@                      @      *@                      &@             �E@      �?      .@      @                      �?                              @              0@               @      �?                      @      *@                      @              ;@      �?      @      @               @      .@      3@              @      $@      �?     �L@      .@     �@@      5@                      @      $@              @      @              (@      @       @      @               @       @      "@                      @      �?     �F@      (@      ?@      ,@              6@     @i@     `p@      ,@      E@      s@     �Q@     �r@      c@     �r@     �i@      :@       @     �]@     �^@      $@      6@     @c@     �A@     @d@     �W@     �d@     @Y@      2@      @     �[@     @[@      $@      3@     `b@      ;@      d@     @S@     `c@     @R@      0@      �?       @      ,@              @      @       @       @      1@      $@      <@       @      ,@     �T@     `a@      @      4@     �b@     �A@     �`@     �M@     @a@     �Z@       @      ,@     �Q@     �]@      @      2@     �]@      ;@     �U@      C@     �Z@      T@       @              *@      5@      �?       @      ?@       @     �H@      5@      ?@      :@              �?     �W@     0q@      (@      $@     �b@      (@     ��@      E@     �y@     @Y@      @      �?      O@     �g@      @      @     �U@      "@     @}@      1@     �q@     @P@       @              .@     �M@       @              $@      �?     `i@      �?     �Y@      2@                      @      9@                       @      �?     @^@              C@      @                       @      A@       @               @             �T@      �?     @P@      *@              �?     �G@     ``@      �?      @      S@       @     �p@      0@     `f@     �G@       @      �?     �E@     ``@              @     �Q@      @     pp@      $@     @f@      F@       @              @              �?              @       @       @      @      �?      @                      @@     @U@      "@      @      O@      @     �d@      9@     @`@      B@      �?              <@     �T@      @      @      L@       @     �c@      5@     �_@      A@                      8@     �R@      @      @     �F@       @      b@      4@     �X@      8@                      @      @                      &@              .@      �?      <@      $@                      @      @       @      �?      @      �?      @      @      @       @      �?              �?                      �?      @              @      @                                      @      @       @               @      �?       @              @       @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO�bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@����Q@�	           ��@       	                   �1@<rB�g�@�           ��@                           �?uWh$�u@�           �@                           �?��fg	 @�            0q@������������������������       �8T���@.            �Q@������������������������       ����ۨ�?z            �i@                          �0@D;��X�@�            �v@������������������������       ����̓@C            �[@������������������������       �-�3��@�            p@
                           �?%*�9��@           z@                           @>O��%�@o            �e@������������������������       ��h��@8            �T@������������������������       ���B��] @7             W@                           �?j�l��E@�            @n@������������������������       �)R�����?/            �S@������������������������       ��I���@n            �d@                           �?��`D@	           L�@                           �?�^ɦ��@           H�@                          �?@�����@           P|@������������������������       ��PZ�7F@           p{@������������������������       ���h%vO@             ,@                           �?e�{�:�@�            @x@������������������������       �^"��@�            �h@������������������������       �^2l�zu@y            �g@                           @��+-P�@�           t�@                           @���h<�@�           X�@������������������������       ���hc~�	@�           ��@������������������������       �
>�1~�@�           P�@                           @��|��@(            �Q@������������������������       ����OA@            �F@������������������������       �#R�@�@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �r@     0�@      D@      K@     `}@     @T@     ��@     �m@     @�@     �t@     �B@       @      H@      `@      �?      $@     @W@      @     �{@     �E@     �l@      L@       @       @      2@     �U@              @      H@      �?     0r@      7@     �`@      ?@       @              @     �B@              �?      8@              b@       @      K@      @       @              @      .@                      .@              2@              .@      @                       @      6@              �?      "@             �_@       @     �C@       @       @       @      *@     �H@              @      8@      �?     `b@      5@     @T@      9@                      @      4@              �?      @              H@      @      2@      "@               @      "@      =@              @      1@      �?     �X@      2@     �O@      0@                      >@     �E@      �?      @     �F@      @     �b@      4@     �W@      9@                      0@      3@      �?              :@       @     �L@      @      C@      (@                      ,@      .@                      1@       @      ,@      @      *@      @                       @      @      �?              "@             �E@              9@       @                      ,@      8@              @      3@       @     @W@      0@      L@      *@                              @              �?       @              E@      @      7@      @                      ,@      4@              @      1@       @     �I@      *@     �@@      $@              $@     @o@     Px@     �C@      F@     �w@      S@     @�@     �h@     �@     0q@     �A@      �?     �N@     �^@      @      @     �U@      ,@      p@      C@      g@     @P@      @      �?     �@@      O@              @      J@      @     �b@      8@     �T@     �B@      �?      �?      =@     �N@               @     �I@      @     �b@      8@      T@     �B@      �?              @      �?              @      �?       @                      @                              <@      N@      @      �?      A@       @     �Z@      ,@     �Y@      <@       @              6@     �D@              �?      :@             �C@      @     �D@      3@       @              @      3@      @               @       @      Q@      @     �N@      "@              "@     �g@     �p@     �A@      C@     0r@      O@     �v@     �c@     �v@     @j@      @@      @     @f@     `p@     �@@      C@     �q@      L@     pv@     @a@     Pv@     �i@      ;@      @     @`@     �e@      :@      @@     �f@     �F@     �_@     �Z@     �b@      a@      4@              H@     @V@      @      @     �Y@      &@      m@      @@     �i@     �P@      @       @      &@      @       @               @      @      �?      4@      @      @      @       @      @      @                      @      �?              0@      @      @      @              @       @       @              @      @      �?      @              @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�Jl!8#@�	           ��@       	                    �?�.0��\@l           X�@                           �?���OX@�           ��@                          �3@=���@�             u@������������������������       �e�
�ҥ @�            �q@������������������������       ��Ցf@&             L@                          �0@m
J�\'@�            t@������������������������       �"���?             >@������������������������       �
l�Vd%@�            0r@
                           �?}��|�@�           �@                           �?��lS��@�            �x@������������������������       �b�e3Y�@g            @d@������������������������       �2��!D{	@�            @m@                           �?�y��Z@�           ȇ@������������������������       ��5e��?@             �I@������������������������       ���k�@�           0�@                           @nX-՚/@*           f�@                            �?�6T �	@1           `�@                           �?�U��+5	@�           ��@������������������������       ��u	��@            �h@������������������������       ��ݏ��	@3           �~@                           �?;G�l�@           @�@������������������������       ���n*��@m             f@������������������������       ��`@ݭ>	@           �{@                            �?A��j@�           ؈@                           �?�����@	            {@������������������������       �~T�*l�@�            `i@������������������������       �C��\�@�            �l@                            @�s!�P@�            �v@������������������������       ��YM�t@�            �l@������������������������       �?p��j@Z            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      9@      L@     �}@      Q@     �@     �h@     ��@     �v@      ;@      @     @X@     @o@      "@      5@     �e@      .@     (�@     �R@     �x@     `b@      $@             �B@     @S@               @      C@             �q@      .@      d@      C@                      &@      >@              @      6@             �e@       @      Q@      2@                       @      :@              @      1@              b@      @     �N@      .@                      @      @               @      @              =@      @      @      @                      :@     �G@              @      0@             �[@      @      W@      4@                              "@                       @              *@              @      @                      :@      C@              @      ,@             @X@      @     @V@      1@              @      N@     �e@      "@      *@      a@      .@     �t@     �M@     �m@     @[@      $@      @      ?@     �D@      @      @     @T@      "@      Q@      ?@     �O@     �G@      $@      �?      (@      6@               @      @@      @      B@       @      =@      0@              @      3@      3@      @      @     �H@      @      @@      7@      A@      ?@      $@              =@     �`@      @       @     �K@      @     Pp@      <@      f@      O@                      @      &@               @      (@      @      @      �?       @      $@                      :@     @^@      @      @     �E@      @     �o@      ;@     �e@      J@              .@     �i@     @t@      0@     �A@     �r@     �J@     �w@     �^@      z@     �j@      1@      .@      d@     �i@      (@      =@     `i@      F@     �d@     �Z@      j@     @b@      $@      @     @U@     @Z@      @      3@     @W@      >@     �S@      Q@      ^@     �R@      @              8@      ?@               @      6@      @      C@      @      H@      5@       @      @     �N@     �R@      @      1@     �Q@      ;@      D@     �N@      R@     �J@      @      &@     �R@     �X@      @      $@     �[@      ,@      V@      C@     @V@      R@      @              ,@      B@      �?      @      >@             �D@      @      @@      *@              &@     �N@     �O@      @      @      T@      ,@     �G@      @@     �L@     �M@      @              G@      ^@      @      @     �W@      "@     �j@      1@      j@     �P@      @              <@     @U@               @      D@       @     �]@      &@      Y@     �E@      @              *@     �A@               @      1@      �?     �P@      @     �C@      7@      @              .@      I@                      7@      �?     �I@       @     �N@      4@                      2@     �A@      @      @     �K@      @     @X@      @     @[@      8@      @              .@      <@      @      �?     �B@      @      K@      @     �P@      *@       @              @      @      �?      @      2@       @     �E@      @      E@      &@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJWhhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @� v�a@�	           ��@       	                   �5@�m���@t           0�@                           �?�2|���@�           p�@                            �?�����@�            �x@������������������������       ���<I��@F            �]@������������������������       �[ó�2�@�            `q@                           @�ʭo3�@�           ��@������������������������       ���_@�k@�            �@������������������������       ��+��>3�?             (@
                           @�BZ��	@�           �@                          �;@-����@�            �@������������������������       �cM��!@1            |@������������������������       �(�n��b	@s            �h@                          �:@�u�b��	@           �{@������������������������       �OOb�	H	@�            �q@������������������������       ���R�.	@h            @c@                           @����1@8           Ě@                           �?�s�iT@�           �@                          �4@�vXs
 @�            pv@������������������������       ����`��?�             n@������������������������       �<�� @K            �]@                           @=�Yq+P@           �@������������������������       ��&��@�           ��@������������������������       ���3��b@�             m@                           @��,(�@9           �~@                          �3@H����/@$           �|@������������������������       �^H��Q@p            �e@������������������������       ��;��	�@�            �q@                          �5@2�ha9�@             A@������������������������       ��f���/@             .@������������������������       �`I��@2@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     Ps@     �@      :@     @P@     �}@     @S@     0�@     �k@     ��@     �u@     �D@      (@     �k@     �s@      1@      I@     �s@      P@     @w@     �f@     �w@     �n@     �@@      @     �R@     @c@      @      7@     `c@      :@     Pp@     @R@      k@     �]@      @              8@     �K@              @      F@      @     �_@      ,@     �V@     �A@                       @      5@              @      "@       @      A@      @     �B@      @                      6@      A@                     �A@      @      W@      &@     �J@      <@              @      I@     �X@      @      4@     �[@      5@     �`@     �M@     �_@     �T@      @      @      I@     �X@      @      4@     �[@      4@     �`@     �M@     �^@     �S@       @                                                      �?                      @      @      @       @     @b@     �c@      $@      ;@     �c@      C@     �[@     @[@     �d@     �_@      <@      @     �R@     �V@      @      *@      Y@      7@      V@      J@     �[@      S@      "@      �?      N@     �O@       @       @     �P@      $@     @S@     �A@     �U@     �A@      @      @      .@      ;@      �?      @      A@      *@      &@      1@      7@     �D@      @      @     �Q@     @Q@      @      ,@      M@      .@      7@     �L@      K@      I@      3@              F@     �J@      @      &@      @@      @      $@     �D@     �B@      <@      3@      @      ;@      0@       @      @      :@      "@      *@      0@      1@      6@                     @V@      m@      "@      .@     @d@      *@     ��@     �C@     0|@      Y@       @             �L@     �e@      @      @     �[@      &@     �|@      7@     �s@      O@      @              .@      B@                      .@       @      g@      @     @V@      ,@                      $@      5@                      @             �a@      �?     �L@      @                      @      .@                      $@       @      F@      @      @@      @                      E@      a@      @      @     �W@      "@      q@      3@     `l@      H@      @              @@     �T@      @       @      T@      "@     �g@      3@     �e@      @@      @              $@     �J@              @      .@             �T@             �J@      0@                      @@     �N@      @      $@      J@       @      a@      0@     �`@      C@      @              :@     �L@      @       @     �H@       @     �`@      &@      `@      A@      @              $@      0@              @      5@             @P@      @      H@      @      @              0@     �D@      @      @      <@       @     �Q@       @     @T@      =@                      @      @      �?       @      @              �?      @      @      @       @               @      @               @       @                                      @       @              @      �?      �?              �?              �?      @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ �-WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @O�IiP@�	           ��@       	                   �5@B�7$��@z           d�@                          �3@��z[�M@�           `�@                           �?�sW��@�           ��@������������������������       ��	�<H@�            pq@������������������������       ��E��X�@           |@                            �?�s�r��@�             x@������������������������       ��#���@�            @k@������������������������       �$'Uˊ0@o            �d@
                           �?�J��'	@�           h�@                            �?��qp�i@�            �r@������������������������       ����_��@C            �Z@������������������������       ��^
�F�@�            @h@                           �?�s!� q	@�           p�@������������������������       �b i���@~            �h@������������������������       ��#k�]	@           H�@                          �2@x[��Y�@K           \�@                           @��T��@b           �@                            �?C)aP��?           �x@������������������������       �u��&�b�?5            @T@������������������������       ���x5 @�            �s@                          �0@���w��@a             c@������������������������       �m8D��?             7@������������������������       �o���k�@S            @`@                            @R���{@�           Б@                          �7@ Ѕv�@p           @�@������������������������       �@�k}��@�            �@������������������������       �8@���@�            @r@                           @{�?+@y            �i@������������������������       ��#'�@              K@������������������������       ��J�&@Y            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �r@     X�@      <@      F@     �}@     @W@     8�@     `k@     H�@     0x@      ;@      &@     @j@     pu@      1@     �A@     �t@      R@     0x@      f@     �v@     Pp@      6@       @     �O@      f@      @      .@      a@      7@     �p@     �V@      j@      \@      @       @      C@     �X@      �?      @      U@      *@     �h@     �P@     �`@     @U@      @       @      &@     �H@                     �B@      @     �S@      1@      F@      @@       @              ;@      I@      �?      @     �G@      @     �]@      I@     �V@     �J@      @              9@     �S@      @      &@     �J@      $@     �R@      7@     �R@      ;@       @              2@      F@      �?      @      <@      @     �D@      &@      J@      *@       @              @      A@      @      @      9@      @     �@@      (@      7@      ,@              "@     `b@     �d@      $@      4@      h@     �H@     @]@     �U@      c@     �b@      .@             �F@     �J@       @      @     �F@      @     �H@      (@      I@      A@      @              0@      2@                      0@      �?      8@              8@      @       @              =@     �A@       @      @      =@       @      9@      (@      :@      =@       @      "@     �Y@     @\@       @      1@     �b@      G@      Q@     �R@     �Y@     �\@      &@      �?      &@      9@      �?      @     �E@      @      7@      0@      4@      C@      @       @     �V@      V@      @      $@     @Z@     �C@     �F@      M@     �T@     @S@      @      �?     �V@     �n@      &@      "@     �a@      5@      �@     �E@     �y@     �_@      @              3@     �R@      @      @      7@             �o@      @     @_@      C@      @              &@      M@       @              $@              i@       @     �V@      5@                              "@                      �?              J@       @      ,@      @                      &@     �H@       @              "@             �b@              S@      2@                       @      0@      �?      @      *@              K@       @     �A@      1@      @                      @                       @              "@              �?      @                       @      (@      �?      @      &@             �F@       @      A@      $@      @      �?     �Q@     @e@       @      @     �]@      5@     `t@     �C@      r@      V@       @      �?     �M@     `c@      @      @      W@      2@     0p@     �B@     �l@     @R@      �?             �B@     �]@      @       @     �L@      .@     �h@      (@     �c@     �E@              �?      6@      B@               @     �A@      @     �O@      9@     �R@      >@      �?              (@      .@       @      �?      ;@      @     �P@       @     �M@      .@      �?               @      @                      ,@      @      *@              *@      �?      �?              $@       @       @      �?      *@              K@       @      G@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�%�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�V�lF?@�	           ��@       	                   �<@��$H\�@w           ��@                           �?���oQ@�           ��@                           �?�<��@�           8�@������������������������       �]Ɖ��@            }@������������������������       ���D@e            �b@                           @Z;��@Q           �@������������������������       �=��u�@/           p�@������������������������       ���0��@"           p}@
                          �>@�0m�L	@�            �q@                            �?�MeaSZ@X            �c@������������������������       ���o��@,            �S@������������������������       �{���-@,             T@                            @A��K�	@K            �_@������������������������       ��ލ)7�@*             O@������������������������       ��}���	@!            @P@                          �6@;(T� @0            �@                           @�G�v��@�           P�@                           �?6ә�@�           ��@������������������������       ��\����?�            �m@������������������������       ��7T@�            @x@                           �?�\G�I@a           �@������������������������       ��I���@�            �i@������������������������       ���i�)@�            Pu@                           �?�M1S@A           �~@                          �8@,�-z�%@�            �m@������������������������       �?�[���@I            @`@������������������������       �?ً�[
@H            �Z@                          �=@ᢎЄ�@�            �o@������������������������       ���|�[@�             k@������������������������       ����_@            �C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@      �@      <@      K@     �|@      T@      �@     @m@     ��@     �v@      =@      &@     `j@     �t@      2@      G@     �s@     �N@      z@     `i@     pv@     �o@      9@      "@      e@     Pr@      $@     �B@      q@      G@     �x@      e@     Pu@     �h@      9@      �?     �J@     @V@              @     @Q@      �?     `f@     �A@     �^@      J@      @      �?     �C@     @T@              @      I@      �?      ]@     �@@     �U@      H@      @              ,@       @              @      3@             �O@       @      B@      @               @     �\@     �i@      $@      >@     �i@     �F@      k@     �`@     @k@     @b@      3@      @     �S@     �\@      "@      1@      c@      =@     �b@     �P@      b@      Y@      &@       @     �B@     �V@      �?      *@     �J@      0@     @P@     �P@     �R@      G@       @       @     �E@      B@       @      "@      E@      .@      5@     �A@      2@      L@                      <@      9@       @      @      2@      "@      @      0@      $@     �D@                      .@      "@              �?       @       @      �?      @      @     �A@                      *@      0@       @      @      0@      @      @      $@      @      @               @      .@      &@      @      @      8@      @      0@      3@       @      .@                      &@      �?                      (@      @      @      (@      @      @               @      @      $@      @      @      (@              "@      @       @       @              @     �R@     �n@      $@       @     `b@      3@     @�@      ?@     �x@     �[@      @              C@     �f@      @      @      T@      "@     �@      2@     Pp@     @P@       @              5@     �T@      @              C@      @     pr@      *@     �a@      :@                      @     �B@                      "@             @b@              B@      @                      1@      G@      @              =@      @     �b@      *@     @Z@      4@                      1@     @X@       @      @      E@      @     �j@      @      ^@     �C@       @              @     �C@              �?      2@             @X@              A@       @      �?              $@      M@       @      @      8@      @     �\@      @     �U@      ?@      �?      @      B@     �P@      @      @     �P@      $@     @[@      *@     �`@      G@       @      @      7@     �A@              @      8@       @      L@      @      O@      7@       @      @      .@      2@                      (@      �?     �@@      �?     �A@      $@       @               @      1@              @      (@      �?      7@      @      ;@      *@                      *@      @@      @             �E@       @     �J@      "@     �Q@      7@                      "@      <@       @              =@       @      I@      @     @P@      2@                      @      @      �?              ,@              @       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@��&�`c@�	           ��@       	                     @���^wO@�           p�@                           �?'�S�2�@W           ��@                           @���YT�@>           @������������������������       �.�ND#�@�            �m@������������������������       �8�E�!��?�            Pp@                            �?`Ǡ��E@           ��@������������������������       �sjeά@�           ؄@������������������������       �Ⱥ���@�             k@
                           @��`�@4           �@                           �?C�&�S2@�            �u@������������������������       ��/�)5@U            �`@������������������������       �����sZ@~            �j@                          �3@,X��� @a            �c@������������������������       �*��c���?Q            @a@������������������������       �d��B�@             5@                          �6@$^��6�@"           ��@                           �?C���J@�           ��@                           �?հt,A@�            �q@������������������������       ���w�2@@             [@������������������������       �Y���@|            `f@                            �?��
I�@�            Ps@������������������������       ���Q���@;            �U@������������������������       ��S|�@�            �k@                           �?y ����@�           d�@                           �?�Ou�i�@�            @w@������������������������       ����@0`@|            `h@������������������������       ���!�p�@h             f@                           @Š�Hw	@�           ��@������������������������       �z (��	@�           0�@������������������������       ��O*�,�@�            �w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `t@     �@      ;@      F@     @|@      Z@     P�@     �i@     0�@     �u@     �A@      @     @Z@     `l@      &@      ,@      h@      7@     ��@     �T@     p|@      `@      &@             @T@     �f@      $@      "@      a@      *@     `}@     @P@     `t@     �T@      @              9@     �L@               @      D@             `l@      .@     �\@      .@      �?              .@      A@              �?      8@             @R@       @     �Q@      &@                      $@      7@              �?      0@             @c@      @     �F@      @      �?              L@     �^@      $@      @     @X@      *@     `n@      I@     `j@      Q@      @              H@     @V@      $@      @     �T@      (@     �d@      >@     �d@     �L@      @               @      A@               @      .@      �?     �S@      4@      G@      &@              @      8@     �G@      �?      @      L@      $@     �c@      1@      `@     �F@      @      @      4@     �@@              @      G@       @      V@      1@     �S@     �C@      @      @      "@      1@                      6@      @      B@      @      9@      ,@              @      &@      0@              @      8@      @      J@      *@      K@      9@      @              @      ,@      �?      �?      $@       @     �Q@              I@      @                      @      (@                      "@             �O@             �F@      @                               @      �?      �?      �?       @       @              @      �?              ,@     �k@     �s@      0@      >@     0p@     @T@     Pu@      _@     �w@      k@      8@      @     @R@     �X@      �?       @     @T@      :@     �`@      3@     @Z@      G@      �?              E@     �B@              @      @@      .@     �T@      @      H@      6@                      =@      3@              @      &@       @      0@      �?      *@      *@                      *@      2@                      5@      *@     �P@      @     �A@      "@              @      ?@      O@      �?      @     �H@      &@      J@      ,@     �L@      8@      �?      �?      @      "@              @      .@      @      .@      @      ,@      $@               @      8@     �J@      �?              A@      @     �B@      "@     �E@      ,@      �?      &@     �b@     �k@      .@      6@     @f@     �K@     �i@     @Z@     `q@     `e@      7@              E@     �K@      �?      @     �C@      @     @S@      3@     �W@     �@@      @              ;@     �@@      �?      @      7@      �?      7@      "@      H@      6@      @              .@      6@                      0@       @      K@      $@      G@      &@      �?      &@     �Z@     �d@      ,@      2@     `a@      J@     @`@     �U@      g@     @a@      2@       @     @Q@     �Y@      *@      $@     �Z@     �G@      H@     @R@      U@      Y@      2@      @     �B@     �O@      �?       @     �@@      @     �T@      *@      Y@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO_�ahG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @C��k�f@�	           ��@       	                   �5@�/�-ؾ@{           ��@                           �?��.��A@�           �@                            �?T�%�H@�             w@������������������������       ���U@J            �]@������������������������       ��rU�7@�            `o@                           �?V��7@�           ��@������������������������       ��x�~Ę@8           P~@������������������������       ��`=@�            `m@
                           @ܑ�u��	@�           �@                           �?�
e�ZV	@           \�@������������������������       �����{@�            0r@������������������������       ��?���	@�           ��@                          �8@{�!�T�@G            �[@������������������������       ��L�@�@             A@������������������������       �I(���@/            @S@                          �4@٘�8�h@5           �@                           @5f=��@S           ��@                           @�o��N�@�            �i@������������������������       �s�EZj@p            `e@������������������������       ���~ħ@             B@                           @��܍�E@�           �@������������������������       �+��?F� @"           �{@������������������������       �91��N@�            Pp@                           @W�7���@�           ��@                            @�
��@[           (�@������������������������       �����@!           �|@������������������������       �f�ȗ�@:             W@                           @(�(@�b@�            `i@������������������������       ���G��6@            �g@������������������������       ���h%vO@             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     (�@      :@     �J@     @{@     �S@     (�@     �m@     ��@     �u@     �E@      0@     �j@     �t@      0@      C@     �r@     �O@      w@     �h@     �z@     @n@     �A@       @     @P@     �d@      @      *@     @b@      3@     �m@     @R@     @n@     �Z@      "@              ;@      H@              �?      @@      �?     @\@      ,@     @Z@      =@                      @      9@                      @              9@      @     �G@      @                      7@      7@              �?      :@      �?      V@       @      M@      7@               @      C@     �]@      @      (@     �\@      2@     �_@     �M@      a@     �S@      "@       @      A@      R@      �?      @      W@      *@     @Q@     �C@     �U@     �K@      "@              @      G@       @      @      6@      @     �L@      4@     �I@      7@               @     `b@     `d@      *@      9@     �c@      F@      `@      _@     `g@     �`@      :@      @      b@      a@      (@      9@     �a@     �B@     �\@     �X@     �f@     @`@      3@              C@      G@      �?      @     �C@       @      H@      3@      O@      ;@      @      @     �Z@     �V@      &@      4@      Z@     �A@     �P@      T@      ^@     �Y@      .@      @      @      :@      �?              ,@      @      .@      9@      @      @      @              �?      .@                      @      @      @       @              �?              @       @      &@      �?              &@      @      (@      1@      @      @      @       @      Y@     �k@      $@      .@     �`@      0@     ��@     �D@     @z@     �Y@       @             �I@     �[@      @      @      M@      @     �x@      3@     �j@      F@      �?              8@      B@                      @      @      U@      @     �C@      "@                      2@      8@                      @      @     �R@              A@      "@                      @      (@                                      "@      @      @                              ;@     �R@      @      @     �I@             �s@      .@     �e@     �A@      �?               @      H@      @      �?      9@             `k@      @     �[@      8@                      3@      :@       @      @      :@              X@      "@     @P@      &@      �?       @     �H@     �[@      @       @     �R@      (@     �h@      6@     �i@     �M@      @       @      9@      S@               @     �J@      "@     @d@      0@     �c@     �C@               @      3@     �R@              @     �I@      "@      _@      &@     �_@     �A@                      @       @              @       @              C@      @      @@      @                      8@      A@      @              6@      @      B@      @     �G@      4@      @              4@     �@@       @              6@             �A@      @     �G@      4@      @              @      �?       @                      @      �?      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ?�BQhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?bU�XGG@�	           ��@       	                    �?)Dq=o/	@           ��@                            �?��C;��@�           �@                           @<^�FÆ@z            �g@������������������������       ���UX��@m            �e@������������������������       �Nɱ���@             ,@                          �9@n\�7@!           p|@������������������������       �4�I��@�            0v@������������������������       ��e
	n�@@             Y@
                           �?Ss�� �	@j           ��@                          �5@��"�@�            �q@������������������������       �k��z��@W            �^@������������������������       �������@g             d@                          �9@8���p:
@�           ؄@������������������������       �Z)�	@'           �|@������������������������       �缠3F
@�            �i@                           �?H%��;@�           "�@                            @��ņ�G@�           ��@                          �4@Sg��?�@�           ȃ@������������������������       ��B��t @�            �w@������������������������       ��3�Lz�@�            �o@                           �?K�[���?_            �c@������������������������       �NL"��<�?9            @X@������������������������       �$8�c�?&            �M@                           @X�f�'@�           �@                          �6@!˷���@�             y@������������������������       �D�R��M@�            �o@������������������������       �A8��m@X            �b@                          �7@�J�)@�           ��@������������������������       �㘖���@           ��@������������������������       �5&���l@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      q@     X�@      >@     �L@      |@      V@     D�@      k@     ��@     �v@      8@      5@     �c@      p@      6@      >@     �m@     �F@     �o@      a@     �k@     �g@      2@       @      H@     �X@      "@      .@     �Y@      "@     `a@      G@     �V@     @T@       @              "@      :@              @      A@      @      F@      1@      B@      .@                      @      9@              @      ?@      �?      F@      ,@      A@      ,@                       @      �?                      @       @              @       @      �?               @     �C@     @R@      "@      &@     @Q@      @     �W@      =@      K@     �P@       @      �?      >@     @Q@       @      "@     �K@       @     @U@      2@     �F@      ?@       @      �?      "@      @      �?       @      ,@      @      $@      &@      "@     �A@              3@     @[@     �c@      *@      .@     �`@      B@      ]@     �V@     �`@     �[@      0@              :@     @Q@       @      @     �B@      �?      F@      4@      G@      >@      �?              (@      7@       @      @      $@             �A@      @      0@      *@      �?              ,@      G@              @      ;@      �?      "@      *@      >@      1@              3@     �T@     �V@      &@      "@     @X@     �A@      R@     �Q@     �U@      T@      .@      &@     �K@     �P@      @      @     �T@      0@     �I@     �H@     �O@      E@      *@       @      <@      7@      @      @      ,@      3@      5@      5@      7@      C@       @      @     �\@     �t@       @      ;@     �j@     �E@     ��@     @T@     Ѐ@     �e@      @              B@     �[@      �?      @     �E@      "@     Pv@      *@     `f@      ?@      @              ?@     @Z@      �?       @     �@@      "@     �p@      (@      b@      :@      @              3@      H@               @      ,@              h@      @     �U@      "@       @              (@     �L@      �?              3@      "@     �R@      @      M@      1@       @              @      @              @      $@             �V@      �?     �A@      @                      @      @              @      @              N@              3@      @                       @      @                      @              ?@      �?      0@                      @     �S@     @k@      @      6@     @e@      A@     �z@      Q@     pv@     �a@       @              9@     �K@      @       @     �G@      4@     @U@     �E@     �S@     �B@                      @     �E@      @      @      =@      @      P@      6@      M@      0@                      4@      (@              @      2@      *@      5@      5@      5@      5@              @      K@     `d@      @      ,@     �^@      ,@     �u@      9@     �q@      Z@       @              B@     �_@      @       @     �P@      ,@     0r@      "@     �i@     �L@       @      @      2@      B@      �?      @     �L@             �J@      0@      S@     �G@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJqeFlhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�&	��@�	           ��@       	                   �5@%46^�@           $�@                           @k�����@�           ��@                            �?L�O��@�            �v@������������������������       �9�.��@�             i@������������������������       ��(��@a             d@                           @���=H*�?�            �x@������������������������       �P����?�            �p@������������������������       �~���p�@R             `@
                          �?@�n�B�@,           p}@                            �?�TT�/@           �{@������������������������       ��Ă-�@Y             c@������������������������       ���]g{@�            Pr@������������������������       ��n�7S@             :@                           �?s�T3t@�            �@                           �?����:
@�           8�@                           @gБb�	@�            0w@������������������������       �� ���	
@�            `l@������������������������       ��w�3 @[             b@                           @^�t7�
@�           ؈@������������������������       ��cі��	@�           ��@������������������������       �w��37	@B            �Z@                           @ĸ�d�@�           ȗ@                           �?g�g�@�            �r@������������������������       �5��d�a@H            �]@������������������������       �UV�W�@p            @f@                          �5@�����0@           (�@������������������������       ���3�a@�           x�@������������������������       � ��H�@:           �}@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     �q@     ��@     �D@      P@     �{@     @T@     �@     �k@     @�@     0v@     �C@      �?     @S@     �f@      @      (@     @[@      @     �{@      @@     @p@     �U@      "@              ?@      \@       @      @      L@             �t@      1@     @d@      A@      @              6@     �I@       @      @      C@             @]@      0@      U@      :@       @              (@      ?@       @      @      0@              M@       @      M@      &@       @              $@      4@                      6@             �M@       @      :@      .@                      "@     �N@              @      2@             `j@      �?     �S@       @      @              @     �D@                      *@             @c@      �?     �G@      @                      @      4@              @      @             �L@              ?@      @      @      �?      G@     �Q@      @      @     �J@      @     @]@      .@     �X@      J@      @      �?     �C@     @Q@      @       @     �I@      @      ]@      &@      X@     �H@      @      �?      "@      5@      @      �?      9@      �?      F@       @      :@      .@       @              >@      H@              �?      :@       @      R@      "@     �Q@      A@      �?              @      �?              @       @       @      �?      @       @      @              2@      j@     �y@      A@      J@      u@      S@      �@     �g@     @~@     �p@      >@      2@     @^@     �e@      9@     �@@     �f@      I@     @^@     ``@      a@     �b@      ;@      @     �G@     @Q@      *@      @     �E@      :@      D@      B@      8@     �L@       @      @      9@      E@      "@      @      8@      4@      @@      (@      4@      @@      @              6@      ;@      @              3@      @       @      8@      @      9@      @      ,@     �R@     �Z@      (@      =@      a@      8@     @T@     �W@     @\@     �V@      3@      &@     �P@     �U@      (@      =@     �]@      1@     �Q@     �S@      Z@      U@      $@      @      @      3@                      2@      @      &@      1@      "@      @      "@              V@     �m@      "@      3@     �c@      :@     p|@     �L@     �u@     @^@      @              4@      L@               @     �C@       @      Q@      6@      J@      7@                      @      1@              @      (@      @      ;@      �?     �A@      *@                      ,@     �C@              @      ;@      @     �D@      5@      1@      $@                      Q@     �f@      "@      &@     �]@      2@     0x@     �A@     pr@     �X@      @              3@     �_@      @      @      G@       @     `q@      3@     @h@      I@       @             �H@     �L@      @      @     @R@      $@     @[@      0@     @Y@      H@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�zhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @�a"/d@�	           ��@       	                     �?���4Z�@�           ��@                           �?�_|@�           �@                           �?���s�@�             j@������������������������       �s!� :@>            @[@������������������������       ��p��D=@D             Y@                           �?F�N_6�@+            }@������������������������       �XS���@�            @u@������������������������       �8�Y$�&@R             _@
                           �?�4��!!	@�           ̘@                          �<@S�Q�@           �|@������������������������       ��K�U�{@�            py@������������������������       ���}��@$            �J@                           @�g�nø	@�           ��@������������������������       �߯���	@p           ��@������������������������       ����?��	@^            �b@                          �4@^���H�@           ԙ@                           @9�z��J@8           �@                           �?c��CO@           �z@������������������������       �<V*��!@�            `m@������������������������       ��N�o���?w            @h@                            �?2QW�*@7           @@������������������������       �j���� @�            pp@������������������������       �:��'@�            �m@                           @F��
ڸ@�           ��@                          �8@� Áj@�           ��@������������������������       ��dz��@           P{@������������������������       �n���2@�            �p@������������������������       ���!+�@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        5@      r@     �@      <@      K@     �~@     �W@     �@     �k@      �@     �t@      D@      4@     �j@     �r@      5@     �B@     @v@      T@     0x@     �f@     Px@     @n@     �B@      @     �H@     @S@      @      *@     �^@      :@     �`@      J@     @]@     �P@      (@              1@      9@              @      8@       @      O@      @      J@      *@      @              @      &@              @      1@       @     �A@      @      2@       @                      $@      ,@                      @              ;@              A@      @      @      @      @@      J@      @       @     �X@      8@     �Q@      G@     @P@      K@      "@      @      ;@      >@      @      @      T@      2@     �A@      D@     �I@     �D@      @              @      6@              @      2@      @     �A@      @      ,@      *@       @      1@     `d@     �k@      2@      8@     @m@      K@     �o@     @`@      q@     �e@      9@             �H@      E@              @     �O@      @      _@      5@     �Y@     �F@      @              E@     �B@              @      J@      @     @^@      1@     �X@      >@      @              @      @              @      &@              @      @      @      .@              1@     �\@     @f@      2@      1@     `e@     �I@     ``@     @[@      e@     @`@      6@      "@      Z@     �b@      2@      .@     �b@      F@      ]@     @U@     �c@     �[@      1@       @      $@      =@               @      4@      @      .@      8@      &@      3@      @      �?      S@     @k@      @      1@     �`@      .@     ��@      D@     �y@     �V@      @              ?@     �^@      �?      $@      B@      @     �{@      3@      l@     �C@      �?              (@     @Q@      �?              (@      @     @h@      (@     �[@      0@                      @     �A@                      "@             �Z@      (@     �L@      (@                       @      A@      �?              @      @      V@             �J@      @                      3@      K@              $@      8@              o@      @     �\@      7@      �?              @      >@              @      (@              `@      @      N@      4@                      ,@      8@              @      (@             �]@      @      K@      @      �?      �?     �F@     �W@      @      @      X@      (@     �h@      5@     �g@      J@       @      �?     �C@     �W@      @      @     @V@       @     `h@      3@     �g@      J@       @      �?     �@@     @P@              @     �N@      @     @_@      @     �[@      8@       @              @      >@      @      @      <@      �?     �Q@      .@     �S@      <@                      @                              @      @      �?       @      �?                �t�bub�k     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�Bx                             �?��ք�<@�	           ��@       	                    �?wX%<�@           ��@                          �6@9���#@�           ؃@                           @��M��@           p{@������������������������       ��GKOn�@r            �e@������������������������       ������?�            �p@                           �?\wέZx@y            �h@������������������������       ����8X�@;            �W@������������������������       �O����;@>            �Y@
                          �5@�x�6q�@�           8�@                          �1@:7 `N@�            �x@������������������������       �p}�B��?W            �a@������������������������       �SOGxg@�            �o@                          �<@���@�            �k@������������������������       ���R`�@r             e@������������������������       ��"J$y@"             K@                           !@��#@�           Τ@                            �?tqlNo@v           ��@                           @
IQ]]�@�           ��@������������������������       ��xgŠV@�            �@������������������������       ���J.	@D             \@                           @i��� �@�           �@������������������������       �D�aϲ�@�           P�@������������������������       �
J���@�           @�@������������������������       ��B=��f@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B`	        "@      s@     @�@      =@     �K@      ~@      W@     d�@      g@     H�@      w@     �E@             �U@     @b@      @      &@     �a@      @     �|@     �@@     �p@     �W@      @              @@     �P@      @      "@     �T@      @     `p@      ,@     @[@      I@                      1@     �E@      �?      @     �G@      @     �j@      $@      S@      7@                      @      7@      �?       @      <@      �?      J@       @      <@      6@                      $@      4@              @      3@      @      d@       @      H@      �?                      .@      7@      @      @     �A@       @      I@      @     �@@      ;@                      "@      &@      @      @      9@              @      @      .@      1@                      @      (@                      $@       @     �E@      �?      2@      $@                      K@      T@       @       @     �M@      �?     `h@      3@     `c@      F@      @              A@      I@                      4@             �c@      @     �X@      ;@                       @       @                      "@             �T@       @      ?@      @                      @@      E@                      &@              S@      @     �P@      5@                      4@      >@       @       @     �C@      �?     �B@      *@     �L@      1@      @              0@      9@       @              ;@      �?      >@      @     �I@       @      @              @      @               @      (@              @       @      @      "@      �?      "@     @k@     `w@      6@      F@     0u@     @U@     ��@      c@     �@     @q@     �C@      "@     �j@     `w@      6@      F@     �t@     @S@     ��@     �b@     �@     @q@      B@      �?     �U@      X@      @      @      W@      8@     �`@      P@     �Z@     �V@      .@      �?     �S@     �U@      @      @     �S@      .@     @^@     �I@     @W@      Q@      (@              "@      $@      @              ,@      "@      *@      *@      ,@      7@      @       @      `@     `q@      .@      C@     `n@     �J@     �|@     @U@     @y@      g@      5@       @     �X@     �f@      *@      :@     �g@      I@     �j@      S@      l@     �`@      5@              =@      X@       @      (@      J@      @     �n@      "@     �f@      J@                      @                              @       @              @       @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJM{�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @8*-�B@�	           ��@       	                    �?�|�|�@r           �@                           �?�S�A�C	@�           |�@                           �?�=샌@�           ��@������������������������       �>0��	@v            �i@������������������������       ����j@           �x@                           �?&^4���	@^           �@������������������������       ���:�I�@�            �s@������������������������       �0,��l
@�            �@
                          �4@�jG�.@�           `�@                          �3@%L�0�I@�            �q@������������������������       �c}��@�            �j@������������������������       ���Z�@*            �P@                          �=@R�����@�             u@������������������������       �:��&�@�            s@������������������������       ��8ǅ&@            �@@                           �?�Ӫ��@H           ��@                          �2@������ @^           Ȁ@                           @�~�V�0�?�            �k@������������������������       ��畢@��?U            �_@������������������������       �&�v���?5            �W@                          �8@o��>�e@�            �s@������������������������       ���(ȋ@�            `o@������������������������       ��k1C�?+            �P@                          �5@8n�v@�           ��@                           @���S@�           ��@������������������������       �46��ʯ@l             f@������������������������       ��)���h@P           `�@                           @un񴉻@.           �~@������������������������       ��;�ʏs@2            @R@������������������������       ��#=�%@�             z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �u@     ��@     �E@      H@     `{@     �R@     h�@      h@     h�@     v@     �C@      (@     �n@     �s@      @@      C@     �q@     �J@     �x@      d@     �v@     �o@     �@@      (@      h@     �k@      <@      @@      k@     �B@      m@     �[@     �o@      i@      >@      �?      N@      W@      �?      $@     �U@      "@     �]@     �@@     �^@     �O@       @              5@      6@                      8@             �O@      @      M@      $@       @      �?     �C@     �Q@      �?      $@      O@      "@      L@      ;@      P@     �J@      @      &@     �`@      `@      ;@      6@     ``@      <@     �\@     �S@     @`@     @a@      6@              D@     �E@      @      @     �A@      �?     �L@      .@     �P@     �G@       @      &@     @W@     �U@      5@      .@      X@      ;@     �L@     �O@      P@     �V@      4@             �J@      X@      @      @     �P@      0@     �c@     �H@     �\@      K@      @              &@     �K@      @      �?      9@      �?     �V@      6@      G@      ;@                      $@      C@                      (@             �S@      2@     �D@      2@                      �?      1@      @      �?      *@      �?      (@      @      @      "@                      E@     �D@              @     �D@      .@     @Q@      ;@      Q@      ;@      @             �B@      D@              @     �@@      &@     �N@      6@      Q@      :@       @              @      �?                       @      @       @      @              �?      �?      �?     @Y@      k@      &@      $@     `c@      5@     ��@     �@@     �y@     �X@      @              4@      N@       @      �?      @@      @     �p@       @     �_@      .@      @              "@      ,@                      $@              a@              H@              @              @      @                                     �V@              8@                              @      @                      $@              G@              8@              @              &@      G@       @      �?      6@      @     �`@       @     �S@      .@                      &@     �E@       @      �?      1@       @      X@      �?     �P@      (@                              @                      @      @     �B@      �?      *@      @              �?     @T@     �c@      "@      "@     �^@      .@     Px@      ?@      r@     �T@      @              =@     �X@      @      @     �L@      &@      p@      $@     `h@     �A@      �?              *@     �B@                      ,@       @      N@      @      >@      $@      �?              0@      O@      @      @     �E@      @     �h@      @     �d@      9@              �?      J@      M@      @      @     �P@      @     �`@      5@     @W@      H@       @      �?      @       @      �?      @      &@       @      2@      $@       @      @                      H@      I@      @      @     �K@       @     �\@      &@     @U@     �D@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJql hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��Jy�Q@�	           ��@       	                   �=@Jifq��@           ��@                           �?+�W�G@�           Ē@                           �?�f�Z�)@�           ��@������������������������       ���Z�@�            @l@������������������������       �*�i�@�            �y@                           �?�mH�n@c           ��@������������������������       �*IH�/�@�            �o@������������������������       ��m�I�@�            `s@
                          �>@:!���@!            �K@������������������������       �\<����@	             (@                           �?���@            �E@������������������������       ���m�`�@             .@������������������������       �9	"�q@             <@                          �3@�a�O6.@�           ¤@                          �1@gI�e�@           `�@                          �0@nMp@�            �u@������������������������       ��S"�_�@J            �[@������������������������       �;�~�5�@�            �m@                           �?������@0           �~@������������������������       ��nr�$�@p             g@������������������������       ��K6�L�@�            `s@                           @�����@u           T�@                          �<@�L�>c�	@�           D�@������������������������       �lg�lc�	@U            �@������������������������       �瑒�X	@q             f@                           @�E�+�@�            �@������������������������       �Yd#��@�           ��@������������������������       �Pu�x�{@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        *@     �q@     `@      :@     �L@     0}@     �S@     ��@      o@     p�@     �w@      B@             @U@     `c@      �?      (@     �_@      @     �z@     �F@     pr@      X@       @             �T@     �b@      �?      @      ]@      @     pz@      A@     Pr@     @T@      @             �B@      R@      �?      @     �N@      @     �o@      5@      `@      J@       @              9@      <@      �?      @      =@      �?      K@      .@      D@      <@       @              (@      F@              @      @@       @     �h@      @      V@      8@                      G@     �S@                     �K@      @     `e@      *@     �d@      =@      @              8@      G@                      C@              H@      $@     @P@      4@      @              6@      @@                      1@      @     �^@      @      Y@      "@      �?               @      @              @      $@      �?      @      &@       @      .@      �?                      @                      �?               @      �?              @      �?               @       @              @      "@      �?      �?      $@       @      &@                                              @      @      �?              @              @                       @       @              �?      @              �?      @       @      @              *@      i@     �u@      9@     �F@     Pu@      R@     0�@     �i@     8�@     �q@      <@      �?      F@     @\@      "@      @     @Q@      (@     @p@     �I@     �g@     �U@      @      �?      2@      F@      �?      @      4@      �?     �`@      5@     �S@      ;@                      "@      ,@               @       @             �G@      @      3@      "@              �?      "@      >@      �?      �?      (@      �?      V@      2@      N@      2@                      :@     @Q@       @       @     �H@      &@     @_@      >@      \@     �M@      @              0@      5@      @      �?      4@      @      ?@      1@      >@     �@@      @              $@      H@      @      �?      =@      @     �W@      *@     �T@      :@              (@     �c@     @m@      0@      D@      q@      N@      t@      c@     �t@     `h@      9@      (@     �^@     @c@      .@     �@@     �g@      G@     �[@      ^@     �c@      _@      2@      @      Y@     �`@      .@      <@     �c@      C@     �X@     @X@      b@      W@      .@      @      7@      3@              @      @@       @      (@      7@      ,@      @@      @             �@@      T@      �?      @     �T@      ,@     `j@     �@@      e@     �Q@      @              ;@      T@      �?      @     @S@      "@      j@      ?@      e@     �Q@      @              @                              @      @       @       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ,�VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @E�T\�:@�	           ��@       	                   �5@"!���@X           ��@                          �1@����K@�           �@                            �?:M?��@�            p@������������������������       ��\�m*@.             S@������������������������       ��S7�al@x            �f@                           �?X�ե��@           �@������������������������       �WB�Q@n           ��@������������������������       �����@�            �m@
                          �:@߾��	@�           ��@                           @������@�           Є@������������������������       ���f�@�            �x@������������������������       ��f�R�		@�            �p@                            �?T��
@           �y@������������������������       ��gj��,	@M            @^@������������������������       ���*�	@�            Pr@                           �?Tܵ٠@@           4�@                          �4@.LÆN� @n           ��@                           @�70�G�?�            �u@������������������������       �A��y�?�            `o@������������������������       ���$�H@B            �W@                          �5@��4Z�@�             k@������������������������       ���r��w�?"             K@������������������������       ��j���@n            `d@                          �8@����;@�           h�@                          �2@����e0@A           ��@������������������������       ���;jL�@�            Pt@������������������������       ���E�@v           ��@                            �?!b\�ml@�            �l@������������������������       �?Q=1�@            �H@������������������������       ��b�[�@u            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      r@     �@      <@      M@     �{@      U@     L�@     �k@      �@     �u@      >@      3@     �i@     u@      7@      C@     �r@      N@     �x@     @e@     pv@      n@      8@       @     @S@     �b@      "@      "@     `c@      1@     pp@     �R@     �j@     �[@      @              &@      C@      �?              =@      �?     �T@      ,@      H@      @@                              0@                       @      �?     �@@       @      ,@       @                      &@      6@      �?              ;@              I@      (@      A@      8@               @     �P@     �[@       @      "@     �_@      0@     �f@     �N@     �d@     �S@      @       @     �J@     �S@      @      @     �W@      (@      ]@     �H@     @[@     �N@      @              *@      @@      �?      @      ?@      @      P@      (@      M@      1@              &@      `@     �g@      ,@      =@      b@     �E@     �`@     �W@      b@     ``@      3@       @     @T@      a@       @      2@     @W@      2@     @X@      J@     �V@     �L@      *@       @     �F@     @S@      @      (@      P@      @     @Q@      .@      Q@      @@       @              B@      N@       @      @      =@      &@      <@     �B@      6@      9@      &@      "@      H@     �I@      @      &@      J@      9@     �A@     �E@      K@     �R@      @              @      1@       @      �?      6@      *@      (@      ,@      1@      ,@      @      "@      F@      A@      @      $@      >@      (@      7@      =@     �B@      N@      �?              U@      j@      @      4@     �a@      8@     @�@     �I@     �{@     @[@      @              *@     @P@              �?      ?@      @     �q@      (@     �_@      8@      �?              &@      <@              �?      *@             �h@      @     �R@      *@      �?              "@      2@                      @             �c@      @      J@       @                       @      $@              �?       @             �E@      @      6@      @      �?               @     �B@                      2@      @     �T@      @     �J@      &@                      �?      1@                      �?      @      :@              @                              �?      4@                      1@      @     �L@      @      H@      &@                     �Q@      b@      @      3@     @[@      1@     �v@     �C@     �s@     @U@      @             �H@     @_@      @      @     �S@      .@     �t@      2@     @p@     �M@      @              ,@     �A@       @      @      .@      �?     �b@      @     �T@      3@                     �A@     �V@       @      @      P@      ,@     @f@      .@      f@      D@      @              6@      3@      �?      (@      >@       @      C@      5@      M@      :@                      �?      @                       @              (@      @      2@      @                      5@      ,@      �?      (@      <@       @      :@      ,@      D@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ8�,IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@%J�R�g@�	           ��@       	                    @�OH�Y4@�           (�@                            �?�w�]@@           �@                           �?
�c R�@�            �q@������������������������       ���\��f@C            �Y@������������������������       ��B����@q            �f@                           �?��|ƻ@�           0�@������������������������       �|����@�             j@������������������������       �_�=�@           `y@
                           @0�{��@B           @�@                           �?���W@�            �k@������������������������       ���(6�@A            @Z@������������������������       ���N��.@I            �\@                           @��FPZ� @�           `�@������������������������       � ��@��?           P|@������������������������       ����TF@�            �l@                           �?�v��Ө@8           ~�@                           �?U����	@z           p�@                            �?�|��@�            �p@������������������������       �_+����@^            �b@������������������������       �UԂ�"@M            �]@                          �:@�`�?
@�           �@������������������������       �8�%���	@<           �@������������������������       �C���X	@�             l@                           @��a���@�           D�@                           �?)�N�'�@�            �s@������������������������       ��9D��@R            �]@������������������������       ����@z             i@                           @Y�%��@�           ��@������������������������       ��Y���@�           ȇ@������������������������       �����@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �r@     0�@      <@      L@     �{@     �U@     Ў@     �m@     Љ@     �u@      =@      "@      Y@      p@      @      1@     �d@      2@     x�@     �S@     pw@      c@      @      "@      Q@     �a@      @      &@     @\@       @      i@     @P@      e@     �Z@      @              8@      J@              �?      =@              N@      8@      Q@      8@       @              @      3@              �?      .@              8@      &@      6@      @                      1@     �@@                      ,@              B@      *@      G@      4@       @      "@      F@     @V@      @      $@      U@       @     �a@     �D@     @Y@     �T@       @              ,@      5@              �?      ?@      �?     �P@      @     �D@      9@      �?      "@      >@      Q@      @      "@     �J@      @     @R@     �A@      N@      M@      �?              @@     �\@              @     �J@      $@     pz@      *@     �i@      G@                      *@     �F@                      $@      @     @V@      @      D@      $@                      @      0@                       @              C@      @      8@      @                      @      =@                       @      @     �I@              0@      @                      3@     �Q@              @     �E@      @     �t@      @     �d@      B@                       @      F@               @      6@             �m@      @     �\@      5@                      &@      :@              @      5@      @      X@      @      J@      .@              .@     �h@     `r@      9@     �C@     @q@      Q@     �v@      d@     0|@     �h@      9@      *@     �]@      c@      1@      8@     �a@      @@     �\@     �[@     �b@     �\@      4@      �?     �D@     �A@       @      @     �B@       @     �E@      0@      L@      7@      @      �?     �@@      ,@      �?       @      3@       @      2@      �?      C@      .@      @               @      5@      �?      @      2@              9@      .@      2@       @              (@     @S@     @]@      .@      1@     �Z@      >@     �Q@     �W@      W@     �V@      0@       @     �J@      V@       @      ,@     @S@      5@      K@      N@     �S@     �D@      (@      @      8@      =@      @      @      =@      "@      1@     �A@      ,@      I@      @       @      T@     �a@       @      .@     �`@      B@      o@      I@     �r@     �T@      @              D@      D@              "@      D@      .@      O@      3@     �O@      >@                      ,@      @              @      .@      @     �@@      @      :@      ,@                      :@     �A@              @      9@      (@      =@      ,@     �B@      0@               @      D@     �Y@       @      @     @W@      5@     `g@      ?@      n@      J@      @       @     �@@     @Y@      @      @     �U@      3@     @g@      :@      n@      J@      @              @      �?      @              @       @      �?      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @|M�9A@�	           ��@       	                   �6@c��ׯ�@x           �@                           �?W���@-           ȓ@                            �?�����@           0z@������������������������       �� iԓ�@�            �n@������������������������       �!�A�y@n            �e@                           �?�7��I�@           x�@������������������������       ��0k�W@�            �q@������������������������       ���mV/�@d           ��@
                           �?�NZ�ڄ	@K           x�@                           �?I�Q1$@�            @m@������������������������       ���(�b@)            �P@������������������������       ����=@k            �d@                           �?عlm,�	@�           (�@������������������������       ���{��@s            @g@������������������������       ����T��	@D           �~@                          �1@'����-@>            �@                           @I�_�?�            �v@                           @��I�%�?�            �q@������������������������       �ޥyx�J�?;            �S@������������������������       ���p/!�?�            �i@                          �0@���@3            �S@������������������������       ��I��ƅ�?             6@������������������������       ��c��MC@&             L@                            @.a��	@O           |�@                           @�m�4g@�           ��@������������������������       �T����@�           H�@������������������������       �3�����@             6@                           @�B�Y%�@�            �n@������������������������       �����' @O            @^@������������������������       �T$���@C            �_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      9@     �M@     0{@      V@     8�@     `j@     Ȉ@     �u@      ?@      4@     `k@     Pt@      1@      F@     r@      P@     0y@     �e@     �v@      n@      6@      &@     �Y@      g@      &@      3@     @c@      3@     s@     �Y@     @m@     @]@      @              8@      L@      �?      @      B@       @     �a@      4@     �X@     �@@      �?              0@      <@      �?      @      1@             @U@      @     @R@      0@      �?               @      <@               @      3@       @     �L@      *@      :@      1@              &@     �S@      `@      $@      ,@     �]@      1@     `d@     �T@     �`@      U@      @      @      9@     �L@      @      @     �E@      "@      J@      2@     �B@      =@               @     �J@      R@      @      $@     �R@       @     �[@      P@     �X@     �K@      @      "@     @]@     �a@      @      9@     �`@     �F@     �X@     �Q@     �_@      _@      .@              5@      >@              @      C@      @     �F@      .@      D@      =@      @              (@      "@                      *@              (@              (@      @       @              "@      5@              @      9@      @     �@@      .@      <@      6@      @      "@      X@     �[@      @      6@     @X@      C@     �J@     �K@     �U@     �W@      "@              9@     �A@       @      @      9@      @      ;@      $@     �@@      2@              "@     �Q@     �R@      @      .@      R@      A@      :@     �F@      K@     @S@      "@              T@     �m@       @      .@     @b@      8@     ؃@     �C@      {@     @[@      "@               @      F@              @      .@             �g@             @U@      ,@       @              @      A@                      $@              d@             �O@      "@                      �?      $@                                      I@              &@      @                      @      8@                      $@             �[@              J@       @                       @      $@              @      @              =@              6@      @       @                      @                                      "@              @      @                       @      @              @      @              4@              2@               @              R@     `h@       @      (@     ``@      8@     �{@     �C@     �u@     �W@      @             @P@     �f@      @       @      \@      4@      v@      C@     �p@     @R@      @             �L@     �f@      @       @     @[@      .@      v@      B@     �p@     @R@      @               @                              @      @       @       @       @                              @      *@      @      @      3@      @     �V@      �?     �S@      6@      @              @      @                       @      �?     �G@             �H@       @      @              @      @      @      @      &@      @      F@      �?      =@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ`^ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��+7�@�	           ��@       	                    �?�j��@           Ȓ@                          �<@���@@7           �}@                           �?2ݭ)@           0z@������������������������       �|�A���@n            �e@������������������������       ��FD�9�@�            �n@                          �=@�-5�٨@#            �J@������������������������       �H�j	"@             :@������������������������       �$��s�@             ;@
                            @i��þ�@�           І@                          �8@LO���&@�           Ђ@������������������������       ��!�L@I            �@������������������������       ���>��@8            �V@                           @�ךf���?U             `@������������������������       �P���� @             C@������������������������       ��<Ս��?<            �V@                           @�n�l@�           .�@                           �?�h{t	@�           ��@                           @����	@�           ̑@������������������������       ����.�	@�           `�@������������������������       �G��@             ;@                            @��ݞ�@           0{@������������������������       ��zUv�@�            �r@������������������������       ���3�Y@P            �`@                           !@C��-�@�           đ@                           @s�JzP@�           ��@������������������������       �ۤ�Z��@�           ��@������������������������       ���W��@�             u@������������������������       ����p���?             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@      t@      �@      =@     �P@     0|@      V@     �@      k@     (�@     �w@     �C@      �?      R@     `e@      @      "@     @Y@      *@      z@     �F@     �p@     �W@      @      �?      I@     �R@      @      @     �J@      @     @X@      >@      X@     �K@       @      �?     �E@     �P@      @      @     �H@      @     @W@      :@      V@     �B@       @      �?      0@      4@                      5@             �I@      @     �E@      0@      �?              ;@     �G@      @      @      <@      @      E@      5@     �F@      5@      �?              @       @                      @              @      @       @      2@                      @       @                       @                       @       @      (@                      �?      @                       @              @       @      @      @                      6@      X@       @      @      H@      @     �s@      .@     �e@     �C@      @              2@      W@       @      @     �B@      @     @o@      ,@     @a@      B@      @              2@      S@       @      @     �@@       @      m@      "@      [@      9@       @                      0@                      @      @      1@      @      >@      &@       @              @      @              �?      &@             @Q@      �?     �A@      @                       @      �?                      "@              0@      �?      "@                               @      @              �?       @             �J@              :@      @              1@      o@     �w@      8@     �L@     �u@     �R@     �@     `e@     �@     �q@     �@@      0@     �f@     @l@      ,@     �A@      p@      N@      k@      a@     �j@      h@      =@      0@      b@      c@      (@      9@     �g@      I@      `@     �X@     �a@     �b@      =@      .@     �a@      c@      (@      9@      g@      I@      `@     �W@     �a@     �b@      5@      �?      @                              @                      @      @      �?       @              B@     @R@       @      $@     @P@      $@      V@      C@     �Q@      E@                      ;@      B@      �?      $@     �K@       @     �I@      :@     �M@      =@                      "@     �B@      �?              $@       @     �B@      (@      (@      *@              �?      Q@     �b@      $@      6@     �W@      .@     Pv@     �A@      r@     �V@      @      �?      Q@     �b@      $@      6@     @W@       @     Pv@     �A@      r@     �V@      @      �?     �D@     @[@      @      @     �K@      @     Pr@      3@     �h@     �K@      @              ;@     �C@      @      0@      C@      @      P@      0@     �V@     �A@      �?                      @                      �?      @                       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ(l-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?nޏ�m@�	           ��@       	                     @����Q@           p�@                          �7@�����Z@K           Ќ@                           �?����4�@�           8�@������������������������       ��e�g�@n             e@������������������������       ��A
&�r @D           �@                           �?���@�            `n@������������������������       �ڡ�Ѓ�@G            �]@������������������������       ��?Yvs�@R            @_@
                          �9@DŧF`�@�             t@                           �?�#�ʮ@�            �p@������������������������       �!��� �@[            �a@������������������������       ������@Q             `@                           @���Z1@%            �J@������������������������       ���`)@             E@������������������������       ���0r��?             &@                           @��c�c@�           ڤ@                           @A�{�r@�           ^�@                           @�G��0	@g           ��@������������������������       �����U
@�            �t@������������������������       �Ƣ��ʤ@�           h�@                          �7@5�>\D�@z           P�@������������������������       �U�,\�@�           ��@������������������������       ��a�@�            @n@                          �3@hG�� �	@�            �s@                           @�`���@0             S@������������������������       �����@#             L@������������������������       �=w�Z�@             4@                           �?:���/�	@�            @n@������������������������       �'h�H	@L            @\@������������������������       �ٶ����@U             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     0r@     ��@      >@      M@     �{@      U@     �@     @m@     H�@     �t@     �D@             �V@     `d@      @      (@     @Y@      (@     @~@      A@     �p@     �P@      "@             @P@      `@      @      @     @R@      (@      v@      6@     @i@      G@      "@             �J@      T@      @       @      I@      @      s@      *@     `a@      7@       @              7@      ;@      @       @      9@      �?     �A@       @     �@@      &@      �?              >@     �J@       @              9@      @     �p@      @     �Z@      (@      �?              (@      H@              @      7@      @      H@      "@     �O@      7@      @              $@      9@              @      *@      �?      (@      @      8@      1@      @               @      7@                      $@      @      B@      @     �C@      @      �?              :@     �A@              @      <@             @`@      (@     @P@      4@                      7@      @@               @      (@             �]@      $@      K@      1@                      .@      0@               @       @             �L@      @      :@      &@                       @      0@                      @              O@      @      <@      @                      @      @              @      0@              &@       @      &@      @                      @      @              @      0@              @       @      @      @                                                                      @              @                      6@      i@     Py@      9@      G@     �u@      R@     �@      i@     �@     �p@      @@      *@     �d@     @v@      5@      G@     Ps@     �K@     p~@     �d@     �}@     �m@      6@      (@     �]@     �k@      0@      <@     @l@     �F@     @g@     @a@     �i@     `d@      4@       @      A@     �G@      @      @      I@      2@     �D@     �C@      A@     �C@      $@      @     @U@     �e@      (@      5@      f@      ;@      b@     �X@     �e@      _@      $@      �?     �G@     �`@      @      2@     �T@      $@     �r@      <@     �p@     @R@       @              <@     �\@      @      *@     �I@      @     �o@      (@     �h@      G@       @      �?      3@      4@      �?      @      @@      @     �H@      0@     @Q@      ;@              "@      A@     �H@      @              B@      1@      N@      A@      B@      =@      $@       @      @      "@                      @       @      ;@       @      ,@       @      �?              @      @                      @       @      8@       @      "@      @               @              @                       @              @              @       @      �?      @      =@      D@      @              >@      .@     �@@      @@      6@      5@      "@      @      "@      .@      �?              4@      @      *@      5@      @      *@      @              4@      9@      @              $@      $@      4@      &@      3@       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�4/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@@ԙ6�S@�	           ��@       	                    �?d��1Sd@W           0�@                          �3@6&�3#�@�           T�@                           �?8�@�@(           �}@������������������������       ������@r            �f@������������������������       �l�**��@�            @r@                           �?nH.��@�           ��@������������������������       �մc���@k            `g@������������������������       �<�B;߁	@           |@
                          �1@��ռ�@�           �@                            �?t_�H� @           p}@������������������������       ��0O����?C             ]@������������������������       ��TC��@�            0v@                           @N�BN)�@�           ��@������������������������       ��D�k�@�           ��@������������������������       �����D;@           Ј@                           @��^!��@A           ��@                           @-��C�@�           �@                           @���=�@R           �@������������������������       ���ެ�-	@�            �w@������������������������       ��:l��@l             e@                           @�}PB�y@�            r@������������������������       �Ag��Ә@L            �^@������������������������       ��5O=9@^            �d@                           �?d��@@E            �[@                           �?&ND�}�@!             K@������������������������       �bE��r @             2@������������������������       �20��C�@             B@                          �;@ENez�@$            �L@������������������������       �0���@            �@@������������������������       ��-9�Dg@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     `r@     x�@      >@     �M@     0}@     �R@     l�@      j@     ��@     �u@      F@      ,@     @j@     �z@      3@      F@     0u@     �D@     ��@     �Y@     Ђ@     �k@      A@      *@     @]@     �c@      (@      8@     �e@      1@      g@      N@      i@     �^@      9@      @     �C@      L@       @      @      Q@      @     �[@     �A@     @R@     �P@      @              (@      @@                      5@             �H@      "@     �A@      7@              @      ;@      8@       @      @     �G@      @     �N@      :@      C@      F@      @      @     �S@     �Y@      $@      3@     �Z@      &@     �R@      9@     �_@      L@      3@              8@     �@@       @       @      2@              A@      @     �L@      @      @      @      K@     @Q@       @      1@     @V@      &@     �D@      2@     �Q@      I@      .@      �?     @W@     �p@      @      4@     �d@      8@     ؆@      E@      y@     �X@      "@              3@      N@              @      8@             �n@      @     �W@      0@       @                      "@              @      @             �T@      �?      (@      @                      3@     �I@               @      4@             @d@      @     �T@      &@       @      �?     �R@     �i@      @      .@     �a@      8@     p~@      B@     0s@     �T@      @      �?      E@     �X@      @      @     @Q@      4@     �d@      9@     @^@      D@      @              @@     @[@      @      "@     �Q@      @      t@      &@     @g@     �E@      @      @      U@     �`@      &@      .@      `@      A@     �`@     �Z@     �c@     @_@      $@      @     �P@      `@      @      .@     @[@      @@     @^@     �T@     �b@      \@      "@      @      D@     �W@      @      @     �R@      ;@     �T@     �G@     �V@     �Q@      @      @      A@     @P@       @      @      M@      6@     �F@      D@     �F@     �I@      @              @      =@      �?      @      0@      @     �B@      @      G@      3@                      ;@      A@      @       @     �A@      @     �C@     �A@      M@      E@       @              0@      .@      @       @      *@      �?      ,@      ,@      ;@      &@                      &@      3@                      6@      @      9@      5@      ?@      ?@       @       @      1@      @      @              3@       @      ,@      8@      "@      *@      �?       @               @       @              "@              "@      1@      @      @      �?                                              @                      @      �?      @      �?       @               @       @              @              "@      &@      @      �?                      1@      @       @              $@       @      @      @      @      @                      (@       @       @                      �?      @      @      @       @                      @       @                      $@      �?              �?      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��!%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Uh$hm^@�	           ��@       	                   �8@�ݥB�p@           ��@                          �4@R�<yO@�           ��@                            �?I{��a@�           ��@������������������������       �����@�            �u@������������������������       ��ᛝ�@�            `s@                           �?�a�F�p@�            `v@������������������������       �&��Ǭ2@{            �g@������������������������       �S%���@h            @e@
                           �?Ź�ͼ�@�            @n@                           �?0Z���@L            @^@������������������������       ���4~@             I@������������������������       ��B�;�@0            �Q@                            @�Y�@G            @^@������������������������       �M����@6             X@������������������������       �j�#0��?             9@                           @E�P]NL@�           ��@                          �9@y(��1	@�           ��@                           @��(~�@�           ��@������������������������       �� �#2�@�           ��@������������������������       ��G$�@
            {@                            �?r	�ʌp	@�            �t@������������������������       �A�� B	@B            �Z@������������������������       ��M0��@�            �k@                          �5@�j�E�@�           ȑ@                          �1@ �x��=@�           @�@������������������������       �;7/6@�            �i@������������������������       ����&@=           �}@                           @#J�{k/@           �|@������������������������       �Y��A=�@�            �r@������������������������       ��ez&��@a            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     pr@     (�@      D@      H@      }@     �U@     ��@     �m@     ��@     �u@      >@             �U@     @f@       @       @     @[@      @     |@      B@     0r@     �S@      @             �P@     @b@       @      �?     �S@      �?     �y@      8@     �k@     �I@      @             �B@     �T@              �?     �H@             r@      3@      b@      ?@      @              :@      I@                      :@             �a@       @     �S@      ,@       @              &@     �@@              �?      7@             @b@      &@     �P@      1@      �?              >@     �O@       @              >@      �?     @^@      @     �S@      4@       @              4@      :@      @              ,@      �?     �R@      �?      D@      @                      $@     �B@      @              0@              G@      @      C@      ,@       @              4@      @@              @      >@      @     �C@      (@      Q@      <@       @              2@      0@              @      5@              (@      @      ;@      ,@                      "@       @                       @              "@              ,@       @                      "@      ,@              @      *@              @      @      *@      @                       @      0@                      "@      @      ;@      @     �D@      ,@       @              �?      0@                       @      @      &@      @     �B@      (@       @              �?                              �?              0@      �?      @       @              *@      j@     0w@      @@      D@     Pv@     @T@     ��@     @i@     ��@     �p@      7@      &@     `a@     `n@      2@      <@     @o@     �M@     �i@     �d@     �j@      e@      3@      @      Z@      g@      1@      7@     �i@     �A@      g@     @]@     �g@      ]@      "@      @     �R@     �Y@      $@      ,@      a@      7@     �^@      J@     @_@     @V@      @       @      >@     �T@      @      "@      Q@      (@     �O@     @P@      P@      ;@      @      @     �A@      M@      �?      @     �F@      8@      3@     �G@      9@     �J@      $@      �?      "@      3@              �?      1@      @      "@      3@      (@      @      @      @      :@     �C@      �?      @      <@      2@      $@      <@      *@      G@      @       @     @Q@      `@      ,@      (@     �Z@      6@     @t@      C@     �s@      Y@      @              6@      T@      @      $@      F@      &@     �l@      6@     �i@      H@       @              @      :@              @      "@             �V@      @     �M@      @                      0@      K@      @      @     �A@      &@     �a@      2@     @b@     �D@       @       @     �G@      H@       @       @     �O@      &@     �W@      0@     @\@      J@       @       @      ?@      ?@      @      �?     �C@       @     �T@      @      S@      9@       @              0@      1@      @      �?      8@      "@      (@      $@     �B@      ;@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�*~hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����H@�	           ��@       	                    �?*��u�@q           F�@                          �<@���:G�@�           0�@                           �?��}���@z           p�@������������������������       �_��)2A@o            �f@������������������������       �Y��!/}@           py@                          �=@>&Yev�@2             V@������������������������       �"S��?             A@������������������������       ���=~�G@             K@
                          �9@���-!D	@�           ��@                           �?L}��i�@�           p�@������������������������       ���>L��@�            @t@������������������������       ���3�@�           ��@                          @A@��#���	@�            z@������������������������       �3R��	@�            �x@������������������������       ��l(�VD@             7@                           @��C���@4           ��@                          �2@T�m�@�           P�@                           @ruY�g�?           @z@������������������������       �̞KO\�?|            `j@������������������������       �dD�����?�             j@                          �9@G*>@�           ��@������������������������       �b��?�@�           P�@������������������������       �������@R            �`@                           �?L�ˍj�@X           ��@                            @�[��jE@~            �i@������������������������       �d�W�Z@^             c@������������������������       ��t��\ @              K@                            @<�����@�            0t@������������������������       �԰x%P@�            �m@������������������������       ��D�gS<@9            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �t@     ��@      >@     �M@     �{@     �T@     ��@     �j@     �@     `w@      1@      2@     �n@     0s@      6@     �F@     �s@      N@     �u@      f@     �x@     pp@      .@      �?      P@     �U@      @      *@     @W@      @     �a@      B@     �c@     �R@      @      �?      L@     �S@      @      &@     �R@      @      a@      :@     `b@      H@      @      �?      1@      ;@                      4@             �H@             �L@      (@                     �C@     �I@      @      &@     �K@      @      V@      :@     �V@      B@      @               @      "@               @      2@              @      $@      $@      :@                      @      @                       @                      �?      @      4@                      @      @               @      0@              @      "@      @      @              1@     �f@     �k@      3@      @@      l@      L@     �i@     �a@     �m@     �g@      &@      $@      _@     �d@      &@      :@      g@      6@     �d@      U@     �h@     �^@      @      �?      8@     �N@      �?      .@     �J@       @      L@      4@      L@      A@      �?      "@      Y@      Z@      $@      &@     ``@      4@     @[@      P@     �a@     @V@      @      @     �L@     �K@       @      @     �D@      A@      D@     �L@     �D@     �P@      @      @     �J@     �H@      @      @      D@      A@      D@     �L@      D@      N@      @      @      @      @       @              �?                              �?      @              �?     �U@     �k@       @      ,@     �_@      7@     ȃ@      B@     p{@     �[@       @      �?     �L@     �c@       @      @     �U@      0@     @~@      1@     pr@      J@      �?              "@     �I@      �?              &@      �?     `l@      @     �X@      1@                       @      >@                      �?      �?     @_@       @     �D@      @                      �?      5@      �?              $@             �Y@      @     �L@      ,@              �?      H@     �Z@      �?      @      S@      .@     p@      (@     �h@     �A@      �?      �?     �B@      W@      �?      �?      M@      &@     �l@      (@     `b@      <@      �?              &@      ,@               @      2@      @      <@              I@      @                      =@     @P@      @      &@      D@      @     �b@      3@      b@     �M@      �?              "@      =@       @       @      (@             �S@      @      J@      2@                      @      :@       @              &@              H@      @      F@      ,@                      @      @               @      �?              ?@      �?       @      @                      4@      B@      @      "@      <@      @     �Q@      .@      W@     �D@      �?              1@      8@      @       @      7@      @      G@      (@     @R@      8@      �?              @      (@      �?      �?      @      �?      8@      @      3@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJP��EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @]Υ�D3@�	           ��@       	                   �3@�����@�           ��@                          �2@�B#��@�           `�@                           @��A56@C           �~@������������������������       ���.��@�             x@������������������������       ���sE�@F            �Y@                           �?��:Y�o@�            `l@������������������������       �Џ�l�v@X            �c@������������������������       ��SQ��@+             Q@
                          �<@�c�\06	@�            �@                           �?���g�@"           ܓ@������������������������       ���E^n@�            �v@������������������������       ��d�;+	@?           P�@                           @�:��	@�            �p@������������������������       ��}D��	@�            @o@������������������������       ����d@             .@                           @�*�;�O@,           ��@                          �2@��u�@�           �@                           �?N�t�\�?           �x@������������������������       ��Al���?�            �i@������������������������       �������?z            �g@                           @�w��:@�           p�@������������������������       ��S�vz@�             r@������������������������       �u����6@.           �|@                           @��>d*[@L           �@                          �=@/�G��@           0y@������������������������       �Dg)ÏW@�            @x@������������������������       �/p3O�@             .@                           @���2�@G             \@������������������������       �RӅ'}@4            �T@������������������������       ���i�*@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �p@     ��@      4@     �K@     �}@     �V@     $�@     `i@     @�@     �v@     �@@      6@     �h@     0t@      &@      F@     �u@     �Q@     �w@      f@     `w@     @q@      <@      @     �@@     �R@      �?      $@     �V@      5@     @g@     �G@     �c@     @V@      @       @      7@     �J@      �?      @     �Q@      @     �a@     �@@     @Z@      G@      @      �?      1@     �A@      �?       @      L@       @     �^@      6@     �W@     �@@              �?      @      2@               @      .@      @      3@      &@      $@      *@      @       @      $@      6@              @      4@      ,@     �F@      ,@     �I@     �E@               @      @       @              @      3@      ,@      ;@      *@      =@      C@                      @      ,@              �?      �?              2@      �?      6@      @              2@     �d@      o@      $@      A@      p@      I@      h@      `@     @k@     `g@      9@      (@     �`@     `j@      @      ;@     �l@     �@@     `f@      X@      h@      `@      5@              :@     �R@              $@     �P@      @      K@      3@      P@     �C@      @      (@     �Z@      a@      @      1@     `d@      ;@     @_@     @S@      `@     �V@      0@      @     �@@     �B@      @      @      <@      1@      ,@     �@@      9@      M@      @      @      @@     �B@      @      @      ;@      ,@      *@      <@      9@      M@       @       @      �?                              �?      @      �?      @                       @      �?      R@     �j@      "@      &@     �_@      4@     p�@      ;@      {@     @V@      @      �?      H@     �b@      @      @     �Q@      *@     P@      *@     `r@     �G@      @              &@     �H@      @              "@             �i@       @     �Y@      ,@                      $@      6@                      @             @Y@       @     �K@      "@                      �?      ;@      @              @             @Z@             �G@      @              �?     �B@     �X@              @      O@      *@     pr@      &@      h@     �@@      @      �?      4@     �E@               @      :@      *@     @V@      @     �Q@      1@      @              1@      L@               @      B@             �i@      @     �^@      0@                      8@     @P@      @      @     �K@      @      c@      ,@     �a@      E@       @              ,@     �M@      @      @      C@      @      `@      ,@     @[@      7@      �?              *@      M@      @      @     �B@      @      `@      ,@     �Z@      1@      �?              �?      �?      @              �?                              @      @                      $@      @              @      1@              8@              ?@      3@      �?              @      @              @      &@              4@              7@      *@                      @                      �?      @              @               @      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�z�'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�yj%�@�	           ��@       	                    �? �,��@�           ��@                           �?�룰`@�           (�@                           �? ����@�            `s@������������������������       ��B�V@�            �k@������������������������       �U4���D@8            �V@                           �?H4���B@�            �v@������������������������       �y����@�            pq@������������������������       ��D5��@5             V@
                           @�\j��<	@�           ��@                          �2@��2�	@x           ĕ@������������������������       ���	�S�@�             r@������������������������       ��[a��h	@�           <�@                          �:@ci��@	@�            `g@������������������������       �<�Y�	�@d             b@������������������������       �rFha�3@            �E@                          �4@f�Pf��@'           ��@                            �?��m^;�@?            �@                          �2@�	Q%1��?�            �k@������������������������       ��&
�\��?R            �]@������������������������       �q���s�?;             Z@                           �?��1�I@�           �@������������������������       ���)����?�            �m@������������������������       �����W�@           0{@                          �7@B�3�%�@�           ��@                          �5@w/wՌ�@�            �v@������������������������       �|0���q@d             c@������������������������       �:�eyr�@�            �j@                           �?��[ُ�@�            �x@������������������������       �u2�,�@s            �f@������������������������       �Oeu�@�            @j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pr@     ��@      1@      L@     �|@      P@     ��@     @m@     8�@     `v@      ?@      5@     �i@     @u@      *@     �C@     �s@     �J@     pz@      h@     Pw@      p@      ;@       @      L@      Z@      �?      "@     @R@      @     �f@      ?@     �b@      O@       @       @      6@     �D@      �?       @      B@       @     @V@      2@      O@      =@               @      1@     �@@      �?      @      ;@       @      J@      0@     �D@      8@                      @       @              @      "@             �B@       @      5@      @                      A@     �O@              �?     �B@      �?     �W@      *@     @V@     �@@       @              9@     �J@              �?      @@              O@      (@      P@      <@       @              "@      $@                      @      �?      @@      �?      9@      @              3@     �b@     �m@      (@      >@     @n@      I@      n@      d@     �k@     @h@      9@      (@     �`@      j@      (@      =@     `j@     �C@     `j@      `@     `j@     �f@      2@       @      3@      F@      �?      �?      @@              U@      :@     �I@      >@              $@     @\@     �d@      &@      <@     `f@     �C@     �_@     �Y@      d@     �b@      2@      @      1@      ;@              �?      ?@      &@      =@      @@      &@      ,@      @       @      .@      7@              �?      9@      &@      6@      6@      &@      @      @      @       @      @                      @              @      $@               @      �?      �?     �V@     `i@      @      1@     �a@      &@     ��@      E@      y@     �Y@      @             �H@     @W@      �?      $@     �K@      @     Pz@      $@     �j@     �B@                      @      4@              �?      $@             �_@       @     �F@      (@                       @      0@              �?      @              R@      �?      0@      @                      @      @                      @              K@      �?      =@      @                     �E@     @R@      �?      "@     �F@      @     pr@       @     @e@      9@                      &@     �@@              @       @             �`@      @      C@       @                      @@      D@      �?      @     �B@      @      d@      @     �`@      1@              �?     �D@     �[@      @      @     �U@      @     @k@      @@     `g@     @P@      @              *@     �O@       @      �?      A@      @      _@      @     �U@      ;@      @                      :@              �?      3@      @      H@      @      B@      "@      @              *@     �B@       @              .@       @      S@       @      I@      2@              �?      <@     �G@      �?      @      J@             �W@      9@     @Y@      C@              �?      .@      7@              @      *@             �I@      (@      J@      *@                      *@      8@      �?      @     �C@             �E@      *@     �H@      9@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ&�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �8@�gB��z@�	           ��@       	                   �3@���V�@b           j�@                           �?����O@�           P�@                           @
}�D@<           @������������������������       ��ZzL @�            �x@������������������������       �|��	@@            @Z@                           @.GL!�@E           �@������������������������       �����v�@�            �v@������������������������       ��3��u@d           ��@
                          �6@�>�S@�           ��@                           @tQ��q_@�           x�@������������������������       ��׭^U�@�           ��@������������������������       �y�փ��@�            �v@                           �?�)�yw@J           �@������������������������       ��JU��@�             k@������������������������       ��~d��F@�            �r@                           �?��)��J	@L           ��@                           �?�/�w�	@;            @                          �?@:�{��@�            @j@������������������������       ���#���@y            �f@������������������������       ��uׅ�d@             <@                           �?F�b �	@�             r@������������������������       ������@4             T@������������������������       �#��&�	@�             j@                           @�`ӆdr@            z@                          �@@�5�= @           �x@������������������������       ��)f�0�@�            �w@������������������������       ��~�.�@	             1@������������������������       �y��-@             6@�t�b�W     h�h5h8K ��h:��R�(KKKK��h��B�
        1@     0s@     ��@      ?@      L@     �}@     �S@     x�@     @k@     ��@     Px@      A@      @     �i@      |@      0@      D@     �u@     �J@     ��@     `a@     X�@      o@      7@      �?     �R@      i@      @      &@     @c@      (@     �|@     �M@     @t@     @\@      $@      �?     �C@      P@      @      "@     �T@      "@     @V@      @@     @V@      Q@      $@              6@      F@      @       @      Q@      @     �S@      7@      U@     �K@              �?      1@      4@      �?      �?      .@       @      &@      "@      @      *@      $@             �A@      a@      @       @     �Q@      @     `w@      ;@     `m@     �F@                      ,@      R@                      ?@      @      ^@      *@      U@      <@                      5@      P@      @       @      D@             �o@      ,@     �b@      1@              @     ``@      o@      "@      =@      h@     �D@     px@      T@     pr@     �`@      *@      @     �T@     �d@      "@      6@     @\@      ?@     �q@     �I@     `i@     �U@      @      @      R@      [@      "@      3@     �U@      :@     �`@      I@     @^@     �I@      @              $@     �L@              @      :@      @     `b@      �?     �T@     �A@              �?     �H@     �T@              @     �S@      $@     @[@      =@      W@     �H@      @              3@      C@              @      H@      @      <@      ,@      >@      9@      @      �?      >@     �F@                      ?@      @     @T@      .@      O@      8@      @      &@     �Y@      _@      .@      0@      `@      :@     @^@     �S@     �a@     �a@      &@      &@      P@      S@      (@      $@     @Q@      ,@     �B@     �J@     �G@     �W@      $@      @      4@      A@      @      @      9@      @       @      7@      5@     �K@       @              1@      @@      @      @      5@      @       @      5@      0@     �I@       @      @      @       @              @      @                       @      @      @              @      F@      E@      @      @      F@      $@      =@      >@      :@      D@       @       @       @      $@      �?              .@       @      .@      @      $@      *@              @      B@      @@      @      @      =@       @      ,@      :@      0@      ;@       @              C@      H@      @      @      N@      (@      U@      :@     �W@      G@      �?              ?@      F@      @      @      L@       @      U@      8@     @W@      G@      �?              :@      F@      @      @      K@      @      U@      5@     �V@      F@      �?              @                               @      @              @       @       @                      @      @                      @      @               @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�[�qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@_�NG��@�	           ��@       	                    @hV,=g@b           R�@                           �?���_�@L           H�@                            �?�&,�}@           �|@������������������������       ���`@O            �_@������������������������       �sp��|�@�            �t@                           @&,�X�@/           0�@������������������������       ��5J�x@t           ��@������������������������       ������@�            s@
                            @�N{f�@           ��@                           �?�jH:�@�           0�@������������������������       ��X���?�            @q@������������������������       ����d�@!            }@                           �?7�c�*@@K            @\@������������������������       ���IM��@+            �Q@������������������������       ���H/E��?             �E@                           �?�z�f@N           ��@                           �?�ҙ^�=	@!            �@                            �?��G~n�@�             q@������������������������       ���"���@9            �U@������������������������       �77M�c@            �g@                          �<@��ԏ	@i           p�@������������������������       ���/��	@           �z@������������������������       ��&?��@R            @`@                           �?��-�r�@-            �@                          �8@��_���@�            �l@������������������������       �fġ��@J            �]@������������������������       �O��&W@L            �[@                           �?7ɜ3@V@�           ؃@������������������������       ����\{@             ?@������������������������       �Wg:��@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@      s@     �@      :@     �F@     `|@      U@     �@     �h@     �@     �v@      4@      @     �`@     �s@       @      7@     @i@      =@     ��@     �U@     @     �f@      @      @     �Z@      k@      @      (@      b@      :@     0u@     �R@     �q@     �a@      @              B@      Q@              @      <@      �?     @b@      1@      ]@     �E@      �?              �?      8@               @      @              A@      @      F@      *@                     �A@      F@               @      7@      �?      \@      ,@      R@      >@      �?      @     �Q@     �b@      @       @      ]@      9@      h@     �L@     �d@     �X@      @      @     �D@      U@      @      @     �T@      2@     �]@      >@     ``@     @S@      @       @      >@     @P@      @      @      A@      @     �R@      ;@      B@      6@      �?              <@     �Y@      �?      &@      M@      @     x@      (@     �j@     �D@                      7@     �X@              "@     �I@             �t@      &@     �f@     �@@                      @      B@               @      0@             �d@      @     �E@      @                      0@      O@              @     �A@             @e@      @     �a@      =@                      @      @      �?       @      @      @     �I@      �?      ?@       @                      @      @      �?       @      @      @      8@              7@      @                      �?      �?                      @              ;@      �?       @       @              @      e@      p@      2@      6@     �o@     �K@     0s@     @\@     �r@     �f@      .@      @      X@     �b@      *@      ,@      a@      ?@     @W@      R@     @Z@     �Y@      *@      �?      9@      M@       @      @      G@      @      I@      3@     �@@      ;@       @              @      *@              @      ,@      �?      2@      &@      0@      @              �?      4@     �F@       @              @@      @      @@       @      1@      7@       @      @     �Q@     @W@      &@      $@     �V@      8@     �E@     �J@      R@     �R@      &@      @     �N@     @Q@      &@      @     @Q@      3@      C@      B@      N@     �F@      $@      �?      $@      8@              @      5@      @      @      1@      (@      >@      �?      �?     @R@     �Z@      @       @      ]@      8@     �j@     �D@     `h@     �S@       @              0@      >@       @              .@      @     �U@      @     �M@      "@      �?              .@      0@       @              @      @      G@              ;@       @                      �?      ,@                       @      @      D@      @      @@      @      �?      �?     �L@     @S@      @       @     @Y@      1@      `@     �B@      a@     @Q@      �?      �?      @       @              @      @      �?              "@      @      @                     �J@     �R@      @      @     @X@      0@      `@      <@     �`@     �P@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@`"pnA@�	           ��@       	                   �1@��җ�@�           ��@                           @��)�n@�           ��@                           �?��'&�@�            u@������������������������       �\T���y@�            pp@������������������������       ��-��R)@+            �R@                            �?C�W��0@�            �r@������������������������       �9��E@n             e@������������������������       ��]b�>@P            ``@
                           @NcB���@           ��@                           @$���b@A           8�@������������������������       �H@��@:           �@������������������������       �������@             .@                           @�|NQ״ @�            �r@������������������������       ��;�@5            �U@������������������������       ��[���r�?�            @j@                           @��K�aD@
           :�@                          �;@�D�4�[	@�           t�@                           �?L����@�           ��@������������������������       ����u	@           |@������������������������       ��ũ��9@�           p�@                          �A@w�a��	@�            �r@������������������������       �U)����	@�            �q@������������������������       ���LЬ1@	             .@                           @��B�<6@f            �@                          �6@췱�:�@�           x�@������������������������       ����Z@�            �t@������������������������       ���;@�!@�            pr@                          �7@�U:��@�            u@������������������������       ��z6�2�@w             g@������������������������       �]��=�@f             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     r@     ��@      >@      F@     �|@     �Q@     ��@      l@     ��@     `w@      @@       @     �R@     �h@      @      @     �`@       @     0@      R@     �t@     �[@      @       @      7@      V@       @      @     �M@             p@      :@      a@      C@                      (@      @@              @      6@             @d@      3@     �P@      5@                      @      ?@              @      3@              `@      &@     �J@      (@                      @      �?                      @             �@@       @      *@      "@               @      &@      L@       @       @     �B@             �W@      @     �Q@      1@               @      @      ?@              �?      5@             �M@      @      =@      ,@                      @      9@       @      �?      0@              B@       @     �D@      @              @      J@     �[@      @       @     �R@       @     @n@      G@     �h@      R@      @      @     �C@     @T@      @      �?     @P@       @      [@     �D@      [@      L@      @      @     �C@     �S@      @      �?     �N@      @      [@     �D@     �Z@      L@      �?      @              @                      @      �?                       @               @              *@      >@              �?      $@             �`@      @      V@      0@                      @      (@                      @              =@      @      >@      @                      @      2@              �?      @             @Z@      �?      M@      *@              0@     �j@     �v@      9@     �B@     Pt@     �O@      �@      c@     `|@     �p@      =@      0@      d@     �n@      4@      =@     �k@     �I@     @j@     �_@      l@     �e@      8@       @      _@     �i@      ,@      :@      f@      B@     �g@     �W@     @h@     �]@      4@      �?      C@      T@      "@      *@      P@      0@      S@      @@      J@     �K@      *@      �?     �U@     �_@      @      *@      \@      4@      \@      O@     �a@     �O@      @      ,@     �B@      C@      @      @     �G@      .@      6@      @@      >@      K@      @      "@     �B@      A@      @      @      F@      .@      6@      @@      <@     �J@      @      @              @                      @                               @      �?                     �J@     @^@      @       @     �Y@      (@      s@      :@     �l@      W@      @              =@     �S@              @     �Q@      @      m@      (@     �a@      G@       @               @      G@               @      D@      @     �`@      @     �Q@      0@       @              5@     �@@               @      ?@             �X@       @      R@      >@                      8@      E@      @      @      ?@      @     �R@      ,@      V@      G@      @               @     �@@      @       @      2@      @     �H@      �?      E@      7@      @              0@      "@       @       @      *@      @      9@      *@      G@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJe��RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@p�gn0@�	           ��@       	                    �?���D�
@|           Ȝ@                            �?\�Sm@�            �@                            �?�	�A�@�             v@������������������������       �Rrkε @j             e@������������������������       �Y�)���@w             g@                          �2@�ڏ��@�            �q@������������������������       ��1@��@u            @h@������������������������       �ɢ>��* @;             W@
                           @�Ӯ��!@�           Ȓ@                            �?�6G�s�@�           `�@������������������������       ��o���@�            �s@������������������������       �q�-�u(@           ؊@                           �?���u@             :@������������������������       ����� � @             (@������������������������       ��|O4l?@             ,@                            @�#�� ~@0           .�@                           @8^T�H@�           $�@                           �?$�t9�r	@�           ��@������������������������       ��a�:�	@n           ��@������������������������       ��  �@�            �j@                           @�ox:��@�           ��@������������������������       �=g�@&           �{@������������������������       �+�>���@~            �g@                           �?:tÒ�@�           p�@                           @��/��@m            �d@������������������������       ���B�\�@S             _@������������������������       ��!��p�?             E@                           @$�ӳ�3	@-           �~@������������������������       ��o[	@            z@������������������������       ��j���@*            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     r@     Ȁ@      <@     �K@     @}@     @S@     �@     �i@     ��@     px@      =@      @     �V@      o@      @      3@      d@      2@     �@      S@     py@     �d@      @              6@     @R@              @     �E@      @     �q@      3@      c@     �C@      �?              0@      F@              �?      ;@             @b@      (@      U@      8@                       @      5@              �?      $@             �R@      @      H@      "@                      ,@      7@                      1@              R@       @      B@      .@                      @      =@              @      0@      @      a@      @     @Q@      .@      �?              @      4@              @      .@       @     @X@      @      C@      @      �?              �?      "@                      �?       @     �C@      �?      ?@       @              @     @Q@      f@      @      .@     �]@      ,@     pv@     �L@     �o@     @_@      @      @     @P@     �e@      @      .@     @\@      ,@     0v@     �L@     �o@      ^@      �?              .@     �D@                      >@      @     �Y@      2@     �R@      ?@      �?      @      I@     �`@      @      .@     �T@      $@     �o@     �C@     @f@     @V@              �?      @      �?                      @              @               @      @      @      �?      @                               @              �?                              @                      �?                      @              @               @      @              &@     �h@      r@      7@      B@     0s@     �M@     `x@      `@     �w@     `l@      7@      @      a@      i@      (@      7@     �h@      E@     Pq@     �U@     0q@     �a@      2@      @      W@     @Y@      "@      1@      \@      A@     �Z@      Q@      a@     @V@      .@      @     �R@     @T@      "@      *@     @V@      4@     �P@      G@     �U@     @Q@      *@              2@      4@              @      7@      ,@     �D@      6@     �H@      4@       @              F@     �X@      @      @     �U@       @     @e@      3@     `a@      K@      @              6@     �Q@       @      @      K@      @     @a@      &@     �X@     �B@                      6@      =@      �?             �@@      @      @@       @      D@      1@      @      @      O@      V@      &@      *@      [@      1@     @\@      E@     @Z@      U@      @              .@      :@      �?      @      4@             �D@      *@      D@      @                      .@      9@      �?      @      2@              ,@      (@      =@      @                              �?                       @              ;@      �?      &@                      @     �G@      O@      $@      $@      V@      1@      R@      =@     @P@     @S@      @      @     �G@      L@      "@      @     �T@      1@     �H@      ;@     �I@     �N@      @                      @      �?      @      @              7@       @      ,@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�$ �E@�	           ��@       	                   �6@�L̤<?@           ,�@                           �?3�>r6�@           ��@                           �?���,�@�            �q@������������������������       ���b�R@P            @_@������������������������       �A�%gF�@d            @d@                           �?Pn�T�� @b           ��@������������������������       �?"P@�            ps@������������������������       �jR�N�3 @�            �o@
                          �<@Y�|�6@�            �w@                            �?-b�@�            �q@������������������������       �-Y�'�@8            @T@������������������������       �tdn�5�@~            @i@                            �?݌�)��@8            @W@������������������������       ���e=�@             ;@������������������������       ��cg.@*            �P@                          �1@F��4;@�           ��@                           @���>*@�            �v@                            �?&��y:@k             f@������������������������       �K�%���@             �H@������������������������       ����i6@K            �_@                            �?,�d @x            �g@������������������������       ��GÁ��?G            @[@������������������������       �+����" @1            �T@                            �?���<��@�           �@                           @���-�}@�           ��@������������������������       ��/!��H@�           (�@������������������������       ��#�A=)@
             1@                          �;@B�Ό!�@*           d�@������������������������       � ��@�           Ԗ@������������������������       �ߔ�߾�	@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     Ps@     �@      ?@     �L@     `{@      T@     �@     �j@     ��@     `u@     �@@             �T@     @e@      @      $@     �X@      @      {@      A@     0s@     �R@      @             �D@      `@      @      @     �N@       @     �u@      *@     �h@     �F@      @              6@      H@      @      @      8@      �?     @T@      &@      Q@      8@       @              @      2@      @              ,@      �?      C@      @      8@      &@       @              .@      >@              @      $@             �E@      @      F@      *@                      3@      T@              @     �B@      �?     �p@       @     ``@      5@      �?              *@      F@              @      :@      �?     �c@      �?      L@      $@                      @      B@                      &@              \@      �?     �R@      &@      �?             �D@      E@      @      @      C@      @     @U@      5@      [@      =@       @              =@      ;@      @      �?      :@       @     @S@      .@     @V@      &@       @               @       @      @      �?      *@      �?      9@      @      .@      �?       @              5@      3@      �?              *@      �?      J@      &@     �R@      $@                      (@      .@               @      (@      �?       @      @      3@      2@                       @      @                       @      �?               @       @      @                      @       @               @      $@               @      @      1@      *@              ,@     `l@     py@      8@     �G@     0u@     �R@     X�@     �f@     H�@     �p@      <@      �?      8@      L@               @      >@              `@      0@     @U@      8@              �?      .@     �@@               @      8@              F@      ,@      <@      .@                      @      @                      �?              *@      @      ,@      @              �?      "@      :@               @      7@              ?@      &@      ,@      $@                      "@      7@                      @             @U@       @     �L@      "@                      �?      $@                      @             �K@       @      =@       @                       @      *@                       @              >@              <@      �?              *@     `i@     �u@      8@     �F@     Ps@     �R@     �z@     �d@     @{@     �n@      <@             �M@      T@      @      $@      V@      4@     �]@     @P@     @\@     �N@      *@             �K@     @S@       @      $@      V@      4@     �]@     �M@     @\@     �N@      $@              @      @      �?                                      @                      @      *@      b@     �p@      5@     �A@     �k@     �K@     @s@      Y@     0t@     �f@      .@      @     �]@     �l@      1@      =@     @h@     �B@      r@     �V@     `r@     �a@      *@      $@      9@      D@      @      @      ;@      2@      2@      "@      =@      D@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�s�"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�E�A@�	           ��@       	                    �?�.	��@           ��@                          �6@�n"D�@*           �@                            �?S�1n@�            `q@������������������������       �J�ґ� @.             R@������������������������       ��\��R@�            �i@                          �;@u:y$�K@{            @l@������������������������       ��8�K�	@U            @c@������������������������       ���3�~@&             R@
                          �>@%#�9��@�           H�@                            @�؈��p@�           ��@������������������������       �{�'��@}           ��@������������������������       �*�.�x�?U            @^@������������������������       ��j��s@             1@                          �5@�R7)&@�           Ф@                          �4@�h;��@�           ��@                           @� `��@�            �@������������������������       �x�u��@�           ؂@������������������������       �EL�G_@_           h�@                           @�	��C@�            �n@������������������������       ��m@!            �N@������������������������       ���2g@t             g@                           @>D&H��@%           ��@                           �?y0X�k�	@           h�@������������������������       �eW���@�            `j@������������������������       ��w-��	@y           Ђ@                          �<@H�_��@$           �{@������������������������       ����r�@�             x@������������������������       ����4!s@*            �M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     pt@     ��@      =@     �G@     �|@     �V@     ��@      j@     ؈@     �u@      5@       @     �S@     �f@               @     �]@      (@     �{@      B@     �q@     �U@      @       @      J@      V@              @     @Q@      @      Z@      9@     @Y@      H@      @              8@      H@              �?      5@      @     @U@      ,@      K@      ;@      �?                      ,@                      @              <@      �?      4@      @                      8@      A@              �?      2@      @     �L@      *@      A@      5@      �?       @      <@      D@              @      H@      �?      3@      &@     �G@      5@      @              1@      =@               @      B@              .@      @      B@       @      @       @      &@      &@              @      (@      �?      @      @      &@      *@                      ;@      W@               @     �H@       @      u@      &@     �f@     �C@      �?              :@      W@               @     �F@      @      u@       @     `f@      @@      �?              9@      V@               @      D@      @     q@      @     @a@      ;@      �?              �?      @                      @             �O@       @     �D@      @                      �?                              @      �?              @      �?      @              1@      o@     �y@      =@     �C@      u@     �S@      �@     �e@     �@      p@      .@      @      W@     `m@      $@      4@     �c@      ?@     @t@      U@     t@     �^@      @      @     �S@     �f@      "@      *@     @`@      3@     @r@     @R@     �o@     @Y@      @      @      I@     �U@      @       @      X@      0@     @X@      O@     @Y@     �Q@      @              <@     �W@      @      @      A@      @     `h@      &@      c@      >@              �?      ,@     �J@      �?      @      :@      (@      @@      &@     �P@      5@      �?              @      (@      �?              (@              "@      @      0@       @              �?      &@     �D@              @      ,@      (@      7@      @     �I@      3@      �?      $@     �c@      f@      3@      3@     �f@     �G@     �k@      V@      h@      a@      &@      $@     �]@      `@      2@      $@     �`@      C@      W@      R@     �U@     @X@      $@      �?      &@      D@              @     �C@      @      A@      0@      <@      @@       @      "@     �Z@      V@      2@      @     �W@     �A@      M@      L@     �M@     @P@       @              C@     �H@      �?      "@     �H@      "@      `@      0@     �Z@     �C@      �?              @@      D@              @     �C@      "@     �^@      0@     @V@      >@      �?              @      "@      �?       @      $@              @              1@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��8<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@{��Nk@�	           ��@       	                    @;����@_           0�@                           �?cz��r@�           ��@                          �1@`���@�            �w@������������������������       ���_n@A            �X@������������������������       ��d� %�@�            �q@                           @�/�e�2@�           x�@������������������������       ��Q���@4           �~@������������������������       ����n�@�             p@
                            �?Mˊ��@�           ��@                           �?r�ˬ^ @�            p@������������������������       ��]��~@P             `@������������������������       �;�[���?G             `@                          �2@[9��Q@           X�@������������������������       �ފ�F@           �z@������������������������       ����@�             x@                          �<@Zqp�E�@=           Ě@                           @�S���t@p           ��@                           @�̲k�@           x�@������������������������       �o���S @~           ��@������������������������       �_�i�T_@�             n@                          �7@s��K�@\           ��@������������������������       �7v��u1@�            �i@������������������������       �q��ڌ@�            Pt@                           @¢
�C	@�             u@                           �?�'��@�            �q@������������������������       ���3@G             ]@������������������������       ��6��s@h             e@                           �?H3!��-@             J@������������������������       �`��� @             ;@������������������������       ���r!w�@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     �~@      :@     �P@     �}@     �U@     ��@     �m@     ��@     �w@      =@      @     @_@     pq@      @      ;@     �m@      C@     h�@     �V@     �~@     �e@      (@      @     �V@     �b@      @      1@     �e@      =@     `p@     @Q@     �j@     �\@       @              A@      F@               @     �B@      @     �]@      .@     �V@      B@                      @      "@                      *@             �H@      @      .@      @                      =@     �A@               @      8@      @     @Q@      (@      S@      @@              @      L@     �Z@      @      .@      a@      9@      b@      K@      _@     �S@       @      @     �@@      N@      @      @     @Y@      3@     @W@      9@      X@     �I@               @      7@      G@      �?       @     �A@      @     �I@      =@      <@      ;@       @             �A@      `@      @      $@     �O@      "@     p|@      5@      q@     �M@      $@              @      =@              @      *@             �a@      @      G@      .@                              ,@              @      "@             �M@      @      8@      .@                      @      .@                      @             @T@      �?      6@                              >@      Y@      @      @      I@      "@     �s@      .@     �l@      F@      $@              &@      F@       @      @      .@      �?      i@       @      ]@      3@      @              3@      L@      �?      @     �A@       @     �\@      @      \@      9@      @      &@     �e@      k@      3@     �C@     �m@     �H@      s@     `b@     pr@     �i@      1@      $@     ``@     �f@      1@      ;@     �g@      =@     0q@     @[@     @p@     �`@      (@      "@     @R@     @Z@      @      1@     @`@      1@      h@     �D@      g@      O@      $@      @     �I@     �U@      @      .@     �T@      (@     �_@      A@     @a@     �D@      $@       @      6@      2@      @       @     �G@      @     �P@      @     �G@      5@              �?      M@     @S@      &@      $@     �N@      (@     �T@      Q@     �R@      R@       @      �?      =@      G@      �?      @      7@      @      :@      5@      ;@      5@      �?              =@      ?@      $@      @      C@      "@     �L@     �G@      H@     �I@      �?      �?      E@      A@       @      (@     �F@      4@      ?@      C@     �A@     �Q@      @      �?     �C@      ?@      �?      $@      B@      2@      *@     �B@      <@     @P@      @      �?      &@      6@               @      3@      (@      @       @      (@      6@                      <@      "@      �?       @      1@      @      @      =@      0@     �E@      @              @      @      �?       @      "@       @      2@      �?      @      @                      �?      @                       @       @      *@              @                               @              �?       @      @              @      �?      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJMw�%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @C$w��(@�	           ��@       	                    �?�U��@y           p�@                           �?�Fb�Y	@�           h�@                            �?nm�~�>@2            ~@������������������������       �ô��R @Y            �a@������������������������       ��_�w	]@�            u@                          �:@�3��2�	@�           �@������������������������       ���8�k	@/           ��@������������������������       �6P�%o	@�            @p@
                          �8@�}�XS�@|           ��@                            �?��r��o@*           p}@������������������������       �<�� �1@Z            `c@������������������������       ��R.�8@�            �s@                           @Sfi�^@R            �`@������������������������       ��|�U>,@G             \@������������������������       ��X�5r� @             7@                           @L\x��@C           D�@                           �?x�UO�@�           x�@                          �4@��N��> @�            px@������������������������       ��Ĳ�o�?�            �p@������������������������       ��(�B��@Q             _@                           @���+��@           ��@������������������������       �B`�q-K@/           �}@������������������������       �`tk��@�            �s@                          �>@��^�v�@D           0@                           �?�u�@9            ~@������������������������       �;���@�             m@������������������������       ���G��@�             o@������������������������       ��(:�"@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     `q@     X�@      >@      P@     0|@      P@     (�@      i@     x�@     �w@      =@      0@     �i@      u@      5@     �I@     �r@      G@     Py@     �d@     @w@     �q@      7@      0@     `d@      n@      3@     �C@      m@     �B@     `o@      `@     Pp@      k@      4@             �K@      R@      �?      @     @R@      �?     �\@      2@      V@      I@       @              2@      8@              �?      .@              D@      @      @@      @       @             �B@      H@      �?      @      M@      �?     �R@      ,@      L@     �E@              0@      [@      e@      2@      A@      d@      B@      a@     �[@     �e@     �d@      2@      $@     �V@     �a@      "@      >@     �`@      5@     �\@     �T@      a@     @Y@      .@      @      2@      ;@      "@      @      :@      .@      5@      =@      B@     �P@      @              F@     @X@       @      (@     @Q@      "@     @c@      C@     �[@     �P@      @              9@     �S@       @      (@     �I@      @     �`@      8@     �V@      H@      @              "@      8@              @      $@       @     �H@      @      ;@      5@      @              0@     �K@       @       @     �D@       @     �T@      2@      P@      ;@                      3@      2@                      2@      @      6@      ,@      4@      3@                      $@      1@                      2@      @      6@      $@      0@      ,@                      "@      �?                                              @      @      @                     �Q@      o@      "@      *@     �b@      2@     ��@      A@     �{@     @X@      @             �F@     `e@      �?      @      Y@      &@      |@      1@      t@     �N@      @              &@     �L@                      6@      @     �h@       @     �T@      ,@                      "@      =@                      &@             �c@              J@      "@                       @      <@                      &@      @      E@       @      >@      @                      A@     �\@      �?      @     �S@      @      o@      .@     �m@     �G@      @              $@     �Q@      �?      @     �G@      @     `b@      $@      c@      8@                      8@      F@                      ?@             �Y@      @     �U@      7@      @              :@     �S@       @      "@     �H@      @      b@      1@     �^@      B@       @              5@      S@      @      "@      H@      @      b@      1@     �^@      =@       @              @      C@      @      @      <@       @      S@      @     �J@      0@                      1@      C@      @       @      4@      @      Q@      *@     @Q@      *@       @              @       @      �?              �?       @                      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ|ǲhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�gmJ�f@�	           ��@       	                    �?��My�>@�           ��@                           @�:(8}n@�           ��@                          �1@/"Sk@�            0s@������������������������       �A��)@8            @X@������������������������       �4s���@            @j@                          �3@��%{��?�            Pv@������������������������       ����3��?�            �q@������������������������       ��e_K8� @)            �Q@
                           �?X�Kidk@�           (�@                           @N�nB.�@           �x@������������������������       �O�����@t            �f@������������������������       ���^�@�            �j@                           @��g:_@�            �@������������������������       �oKF߫]@�            @t@������������������������       �*W0��9@           �{@                            �?��R�Z�@2           N�@                           @
���/�@�           �@                           �?���n�O	@�           X�@������������������������       �EXԏP�@�            �h@������������������������       �?��@_�	@2           p~@                           �?�B�2�@�            �x@������������������������       �KR�p�@R            @_@������������������������       ��r*��l@�             q@                          �<@��Tï@           h�@                          �9@f�(��S@           ��@������������������������       ����,Z�@�           �@������������������������       ��ʠ���@�            �k@                           @JX�n5	@s            �e@������������������������       �oT�T�	@S             `@������������������������       �����@             �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     `r@     �@      ;@     �O@     P}@     �T@     ��@     `o@     x�@     �t@      :@      @      [@      m@      &@      4@     �e@      &@     ��@     @V@      y@     �a@      @             �A@     �V@              @     �F@      �?     �r@      .@      a@     �A@       @              9@     �B@              @     �A@      �?     �V@      ,@      R@      ;@      �?              @      &@                      $@             �F@       @      6@       @                      4@      :@              @      9@      �?      G@      (@      I@      9@      �?              $@     �J@              �?      $@              j@      �?      P@       @      �?              @      D@                      @             �e@      �?      K@      @      �?              @      *@              �?      @             �A@              $@      �?              @     @R@     �a@      &@      .@      `@      $@     �t@     �R@     �p@     @Z@      @      @      @@     �F@      @      @      R@      @      L@     �F@     @R@      G@      @       @      *@      :@      @      @     �@@              B@      @      B@      0@      �?      �?      3@      3@               @     �C@      @      4@      C@     �B@      >@      @             �D@     �X@      @       @     �L@      @      q@      =@     �g@     �M@                      5@     �I@      �?       @      =@      @     �X@      6@     @R@      6@                      4@     �G@      @      @      <@      �?     �e@      @     �]@     �B@              4@     @g@     �s@      0@     �E@     pr@      R@     x@     @d@     �w@     @h@      3@      "@      Z@     �d@      @      4@     �a@      F@      h@     @X@     �i@     �W@      @      "@     �T@     @X@      @      0@      Z@      B@     �T@     @S@     �Z@      P@      @              <@      6@              @      8@      �?     �D@      @      K@      1@              "@     �K@     �R@      @      *@      T@     �A@      E@     �Q@      J@     �G@      @              5@      Q@      @      @      B@       @     @[@      4@     �X@      >@      �?                      0@       @              $@      �?     �C@      @      B@      ,@                      5@      J@       @      @      :@      @     �Q@      *@      O@      0@      �?      &@     �T@     `b@      "@      7@     `c@      <@      h@     @P@     `f@      Y@      *@      @      O@     �_@      @      2@     @]@      4@     �e@      H@     �c@      T@      *@      @     �G@     @X@      @      *@      X@      $@     �`@      ?@     �Z@     �M@      "@      @      .@      =@       @      @      5@      $@     �D@      1@      J@      5@      @      @      4@      5@       @      @      C@       @      3@      1@      4@      4@              @      *@      2@       @      @      :@       @       @      1@      *@      .@                      @      @                      (@              &@              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJbzymhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�6Bk]@�	           ��@       	                   �3@���@X           �@                           @"��@�           �@                           @ka��x@�            �v@������������������������       �V6)S�@�            �r@������������������������       ���䯁�@+            �P@                          �1@��+13 @�            `u@������������������������       ���*�K��?f            @e@������������������������       �Ͻ@6�} @n            �e@
                          @@@��ʡA@�           �@                          �7@�JC��@�           ��@������������������������       �������@f           x�@������������������������       ����9��@.           �@                            @�G �]@             :@������������������������       ��I��,�?             *@������������������������       ��D����@	             *@                           �?b�_��@A           ��@                           �?�dHɞ1	@{           X�@                          �<@P5pq��@�            �p@������������������������       ��A#�).@�             o@������������������������       �C�H�IO@             7@                           �?��d*�	@�           ��@������������������������       ���#��	@�            p@������������������������       ����	@5           �}@                            �?V���b@�           l�@                          �4@��i���@�            �q@������������������������       ��5v� ��?a             a@������������������������       ��~�T�@Y            �b@                          �9@ד��_@           ��@������������������������       ����32@�           h�@������������������������       ���ys@Y             b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@     ��@      5@     �N@     @}@     @X@     ��@     �i@      �@     �v@      ?@       @     �`@     �p@      "@      ;@      i@      F@     �@     �T@     0u@     �d@      *@             �D@     �V@      �?       @      K@      @     �p@      3@     @e@      K@                      <@     �M@                      A@      @     @X@      1@     @T@      E@                      .@      J@                      >@      @     �T@      $@     @R@      ?@                      *@      @                      @      @      ,@      @       @      &@                      *@      @@      �?       @      4@             `e@       @     @V@      (@                      $@      .@               @       @             �U@              G@       @                      @      1@      �?              (@              U@       @     �E@      $@               @     �V@     `f@       @      9@     `b@      C@      n@     �O@      e@     @\@      *@             �V@     �e@       @      7@     @b@      ?@      n@     �O@     �d@     �[@      *@             �E@     @Y@      @      2@      W@      6@     �`@      4@     �T@     �B@      @             �G@      R@       @      @      K@      "@     �Z@     �E@     �T@     �R@      "@       @      �?      @               @      �?      @                      @       @                      �?      @                              @                      �?                       @               @               @      �?                              @       @              ,@      e@     �r@      (@      A@     �p@     �J@     0}@      _@     }@      i@      2@      ,@     @Z@      b@      "@      5@     �d@      =@     �`@     �R@     �e@      ]@      1@              A@     �H@               @      @@              N@      ,@     �L@      7@                      >@      H@                      9@             �M@      ,@     �J@      3@                      @      �?               @      @              �?              @      @              ,@     �Q@      X@      "@      3@     �`@      =@     �R@     �N@     �\@     @W@      1@       @      6@      E@      @      $@      C@      @      ;@      5@      D@     �E@      @      (@     �H@      K@      @      "@     �W@      7@      H@      D@     �R@      I@      ,@             �O@     �b@      @      *@     �Y@      8@     �t@     �H@     Pr@      U@      �?              .@     �C@      �?      @      &@      "@     �Z@      ,@      N@      :@                      @      3@                      @      �?     @S@       @      4@      @                      &@      4@      �?      @      @       @      =@      (@      D@      3@                      H@      \@       @      "@     �V@      .@     @l@     �A@      m@      M@      �?              @@      X@       @      @      M@      @      k@      9@      i@     �E@      �?              0@      0@              @     �@@      "@      $@      $@      @@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJpJ
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?t���F@�	           ��@       	                    �?`e��~@           8�@                          �<@�:��^&@;           �~@                           �?�F��c�@           �{@������������������������       ����ž�@k            �d@������������������������       �̵���@�            `q@                          �?@�(�	�@#             I@������������������������       �J,Gz"�@             E@������������������������       �      �?              @
                           @{l�ԉn@�           ��@                            �?���=� @g           ��@������������������������       �4��( @`            �c@������������������������       ���m�'z @           Py@                          �6@��d#@q            �e@������������������������       ��C"�l�@L             [@������������������������       ��X���� @%            �P@                           @���<�3@�           ��@                            @��ɲh�	@�           `�@                           @�O_(z	@g           �@������������������������       ��9�q�-	@r           �@������������������������       ��y��D	@�            �w@                           �?zBH�	@�           ؂@������������������������       ��U�0�	@>           p~@������������������������       �+7Z�D@I             ]@                          �;@�-qw�@�           ��@                           @�*9�fo@�           d�@������������������������       ���@3           Ќ@������������������������       ��h���@U            �_@                            �?��69��@4            �R@������������������������       ����b��@            �C@������������������������       ���Xl�N@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     q@     ��@      :@     �N@     px@     �U@     L�@     �l@     ��@     �v@     �B@             �T@     `e@      @      "@      T@      ,@     �{@     �E@     r@     @U@      @             �J@     �V@       @      @      G@      @     @X@      @@     �Y@     �L@       @              F@     �T@       @      @     �C@      @     �W@      =@      Y@      D@       @              "@      B@                      ,@              C@      @      J@      *@                     �A@     �G@       @      @      9@      @     �L@      8@      H@      ;@       @              "@      @              @      @               @      @       @      1@                      @      @              �?      @               @      @      �?      1@                      @      �?               @                                      �?                              >@     @T@      @       @      A@      @     �u@      &@     `g@      <@      @              9@      M@              �?      :@      @     �q@      @     �`@      2@      �?               @      4@              �?      @       @     @S@              D@       @      �?              7@      C@                      5@      @      j@      @     �W@      $@                      @      7@      @      �?       @              P@      @     �J@      $@       @              @      ,@              �?       @              H@      �?      7@      @       @                      "@      @                              0@      @      >@      @              6@     �g@     �x@      5@      J@     ps@      R@     ��@     @g@     ��@     pq@      @@      6@     �`@      n@      2@      D@     �k@     �L@     �l@      c@     @n@     �e@      <@      "@     @T@     �_@      $@      >@     �a@      =@     �b@      Z@     `b@     @\@      1@      @      M@     @P@      @      3@      V@      7@     @T@      H@     �Y@     �S@      @      @      7@     �N@      @      &@     �J@      @     @Q@      L@     �F@      A@      (@      *@     �J@     �\@       @      $@     �T@      <@      T@      H@     �W@     �N@      &@      *@     �F@     �T@      @       @     @R@      9@     �L@      B@     �T@      H@      &@               @      ?@       @       @      "@      @      7@      (@      *@      *@                      L@      c@      @      (@      V@      .@     �v@      A@     �q@     @Z@      @             �I@     �`@      @      "@     @Q@      ,@     �v@      @@     0q@     �X@      @             �B@     @^@      �?       @     @P@      &@     �s@      ;@     �o@     �T@       @              ,@      &@       @      �?      @      @      H@      @      5@      0@       @              @      4@              @      3@      �?      @       @      (@      @                      @      .@                       @                      �?       @      @                       @      @              @      &@      �?      @      �?      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�����L@�	           ��@       	                    @&�Cɳ�@           ��@                           �?G�EA�@'           ��@                           �?E��K@1           ��@������������������������       ��[ �@�            @t@������������������������       ��y����@W           Ѐ@                           @�f �Y�@�            �x@������������������������       �2��@�            p@������������������������       �A#s$�w@X            �a@
                           �?�5��aP@�           <�@                            �?`*n�a�?           �{@������������������������       �g�"�`�?E            �X@������������������������       �D ښm @�            �u@                          �4@!�d�@�           ��@������������������������       ��:�%@c           �@������������������������       ���^̶@w             f@                           �?���H		@�           8�@                           �?%�s�`\@�            �w@                          �<@w��[M@s            �f@������������������������       ��Q���`@Y            �`@������������������������       �P���?@             H@                           @GU�Z�h@~            �h@������������������������       �EO��K4@P            @]@������������������������       ���,�N@.            @T@                           @�q���y	@�           L�@                           @�tA��B	@8           ��@������������������������       �J�:Aؿ	@s           ��@������������������������       ��<�Ƽ�@�            �s@                          �8@�T^	@r            @h@������������������������       ���RΔ@*             R@������������������������       �ZSn&��	@H            �^@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     �q@     Ђ@     �A@      M@     `|@     �W@     �@      j@     ��@     �u@      >@      @     @b@     w@      0@      :@     0q@     �E@     Ј@      Y@     �}@     �e@      @      @     �[@     `i@      *@      1@      g@     �A@      r@     �S@     �h@     �_@       @      @      W@      a@       @      .@     �a@      :@     �c@     �L@      `@     @W@       @              5@     �M@      �?      @     �H@      @     �T@      4@      H@      >@              @     �Q@     @S@      @       @      W@      3@      S@     �B@     @T@     �O@       @              3@     �P@      @       @      F@      "@     @`@      5@      Q@     �@@                      0@      ?@               @      <@      @     @W@      "@      F@      =@                      @      B@      @              0@      @     �B@      (@      8@      @                     �A@     �d@      @      "@     �V@       @     �@      6@     pq@     �G@       @              "@      N@              @      4@      �?     �n@      "@     @U@      (@                              3@                      �?             �O@              (@      @                      "@     �D@              @      3@      �?     �f@      "@     @R@      "@                      :@     �Z@      @      @     �Q@      @     `p@      *@     @h@     �A@       @              9@     �S@      �?      @      H@      @     �i@      $@     �a@      >@                      �?      ;@       @       @      6@      @     �K@      @      K@      @       @      @     �a@      m@      3@      @@     `f@      J@     @m@      [@     pq@      f@      :@      �?      ?@     �P@       @      "@      B@      @      Y@      $@      U@     �@@      @      �?      4@     �D@              "@      8@              7@      @      @@      7@       @      �?      2@      :@              @      4@              6@       @      >@      "@       @               @      .@              @      @              �?      @       @      ,@                      &@      :@       @              (@      @     @S@      @      J@      $@      �?              $@      $@                      @      @     �H@      @      =@      @      �?              �?      0@       @              @              <@      �?      7@      @              @     �[@     �d@      1@      7@     �a@     �H@     �`@     �X@     `h@      b@      7@       @      U@     @_@      0@      7@     �]@      D@      \@     �R@     �e@     �`@      *@      �?      Q@      T@      ,@      .@      T@      B@     �E@     �M@      W@     �W@      *@      �?      0@     �F@       @       @     �C@      @     @Q@      0@      T@     �B@              @      :@     �D@      �?              8@      "@      6@      7@      7@      (@      $@              @      =@                      *@      @       @      @       @      @      �?      @      5@      (@      �?              &@      @      ,@      0@      5@      "@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��V4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�XE���@�	           ��@       	                   �;@��y�	@d           <�@                          �1@��5�+�@�           p�@                           @������@�             q@������������������������       �
{r6�]@y            �h@������������������������       �v칒*@.            �R@                           �?�w��l�@�           (�@������������������������       �6I�Z��@+           �}@������������������������       ��5��~	@�           ��@
                            �?l��֠�	@�             t@                          �=@)�}[�`
@:            @W@������������������������       �C�P�V�@            �D@������������������������       �>����-@              J@                            �?qMx
O	@�            �l@������������������������       ��g��@1             T@������������������������       ��$��=	@d            �b@                           @���/@4           ��@                           @��MU@�           X�@                            �?+���l.@�            �x@������������������������       ���託�@F            �Z@������������������������       �F�՗@�@�             r@                           @G�C�@�           P�@������������������������       ����Ш)@*           p~@������������������������       ��T ��@�            0r@                           �?�DϻP @U           ��@                           �?O����+@�             i@������������������������       ���v$B@J            �[@������������������������       �]DW-��@8            �V@                           @�h��@�            �t@������������������������       ��ԝ�$@�            �q@������������������������       �����h	@             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      r@     ȁ@     �B@      P@     0|@     �S@     ؎@      l@     P�@     �w@     �A@      0@     �h@     �s@      ?@     �G@     �t@      L@     �u@     �g@     �w@     `p@      ?@      "@     `c@     @q@      6@      C@     �q@     �E@     �t@      c@     �u@      i@      :@       @      ,@     �C@      @      �?      ?@      �?     @T@      5@      N@      5@                      @      8@      @      �?      5@             @P@      ,@     �J@      &@               @      @      .@                      $@      �?      0@      @      @      $@              @     �a@     �m@      3@     �B@     �o@      E@     �o@     ``@     �q@     �f@      :@              @@     �P@      @      @      I@      @      `@      4@     �^@     �E@              @     @[@     @e@      .@      @@     @i@     �B@     �^@     �[@     �d@      a@      :@      @     �E@     �D@      "@      "@     �F@      *@      1@      B@      B@     �N@      @       @      @      ,@      @      �?      ,@      "@      @      $@      "@      .@      @       @              @      @      �?       @      @      @       @       @       @                      @      $@                      (@      @      @       @      �?      @      @      @      C@      ;@      @       @      ?@      @      $@      :@      ;@      G@       @      �?      ,@      @      �?      @      @               @      1@      *@      2@              @      8@      4@      @      @      <@      @       @      "@      ,@      <@       @       @      W@     �o@      @      1@     �^@      7@     �@      B@     �x@     �]@      @       @     �N@     �f@      @      @     �P@      .@     @~@      1@     �p@     �P@       @       @      :@      T@      @      @      ;@      ,@     �a@      "@      P@      ;@                       @      3@      @              @              H@       @      ,@       @               @      2@     �N@              @      7@      ,@     @W@      @      I@      3@                     �A@      Y@              @      D@      �?     pu@       @     �i@      D@       @              :@      H@                      6@      �?     �l@      @     �^@      <@       @              "@      J@              @      2@             @\@      �?     �T@      (@                      ?@      R@      @      $@      L@       @      c@      3@     �_@      J@       @              @      8@               @      (@      �?      W@       @      H@       @       @              @      1@               @      @      �?      L@      @      4@      @                              @                       @              B@      @      <@      @       @              ;@      H@      @       @      F@      @     �N@      &@     �S@      F@                      4@     �E@              @     �A@      @     �L@       @     �Q@      E@                      @      @      @      @      "@       @      @      @       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�0'*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@(�ُ�@�	           ��@       	                    @X��,/@#           N�@                           �?t�=�@(           ��@                          �3@S��`��@�            Px@������������������������       ����@�            @n@������������������������       ���0r�@\            `b@                           �?�]��	�@)           H�@������������������������       ��0��	@�           (�@������������������������       ����:7�@�            @p@
                           @�/zΦ@�           �@                          �1@� 2�@�            �q@������������������������       ����{;�?1             S@������������������������       �X�.F1@�             j@                           @QO���@J           �@������������������������       �lX��0{ @o           H�@������������������������       �v.m�d@�            @u@                          �<@׹�!Q	@�           ��@                          �7@�ܨ{�@�           �@                           �?�\��@�            �l@������������������������       ��1t��f@B             [@������������������������       �����@O            @^@                           �?��7Y߀@           ��@������������������������       ����ӔH	@�            0{@������������������������       �f�����@           �z@                           @�K�1�	@�            v@                            �?�6���@�            @k@������������������������       �ԥ�Fڷ@M            @^@������������������������       �N�Z�}-@?            @X@                           �?��]m{	@V            �`@������������������������       ���ּ �	@2             S@������������������������       �7����k@$            �M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     Ps@     p�@     �B@      K@     �~@     �S@     Ў@      n@     ��@     �u@      F@      @     `e@     �t@      .@      >@      p@     �@@     h�@     @_@     X�@      g@      ,@      @     �^@     �e@      &@      3@     `f@      8@     p@     �Z@     �m@     �\@      &@              C@     �F@       @       @     �F@      @     �[@      6@     �W@      8@      �?              5@      =@              �?      :@       @     �Q@      @     �O@      7@                      1@      0@       @      �?      3@       @      D@      0@      @@      �?      �?      @     @U@     @`@      "@      1@     �`@      4@     @b@      U@     �a@     �V@      $@      @     @R@     �T@      @      ,@      Y@      &@      U@      I@      Y@     �R@      $@              (@     �G@       @      @      A@      "@      O@      A@      E@      .@                      H@     �c@      @      &@     @S@      "@     `�@      3@     �q@     �Q@      @              3@      K@      �?              0@      @     �[@      @     �J@      0@       @              �?      &@                      @             �F@      �?      &@      @                      2@     �E@      �?              *@      @     @P@      @      E@      (@       @              =@      Z@      @      &@     �N@       @     �y@      *@      m@      K@      �?              0@      M@      �?      @      >@             �q@      @      c@     �A@                      *@      G@       @      @      ?@       @      `@      "@     @T@      3@      �?      @     @a@      h@      6@      8@     �m@     �F@     �i@     �\@     pp@     �d@      >@      @     @X@     �b@      1@      &@     `f@      ?@     �e@      U@     @l@     �X@      7@              >@     �G@      @      @      B@      @      >@       @      D@      6@      @              (@      8@       @      �?      8@      �?      @      @      ,@      0@      @              2@      7@      �?       @      (@      @      9@      @      :@      @      �?      @     �P@     @Y@      ,@       @     �a@      :@     �a@      S@     @g@      S@      2@       @      D@      I@      *@      @     �V@      .@     �E@     �H@     @R@      D@      0@      �?      ;@     �I@      �?      @      J@      &@     �X@      ;@     @\@      B@       @       @     �D@     �F@      @      *@     �L@      ,@     �@@      ?@     �B@      Q@      @      �?      ,@      >@       @      @      D@      &@      5@      0@      5@     �I@      @               @      *@              @      .@      $@      (@      &@      &@      @@      @      �?      @      1@       @       @      9@      �?      "@      @      $@      3@              �?      ;@      .@      @       @      1@      @      (@      .@      0@      1@      �?      �?      *@      "@      @       @      @       @      @      ,@      @      &@      �?              ,@      @                      (@      �?      "@      �?      $@      @        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ ��9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @XSR/E@�	           ��@       	                    @u�*Bb�@�           ��@                          �;@�J7+�@h           Е@                           �?�Q� @�           p�@������������������������       ���W2T@�            `w@������������������������       ��:`�@�           0�@                           @�;��i�@�             k@������������������������       ����q@K            @_@������������������������       �w�J��A@8            �V@
                          �4@�����@j           ��@                           �?q����@�           �@������������������������       ������?�            0s@������������������������       �"�]1 @.            }@                           @L��J��@�            �@������������������������       ��D�FF�@\            `a@������������������������       �l-��@,           P}@                          �3@AS��:�@�           ȑ@                           @"��$�@�            Pw@                           �?�Hď��@�            @o@������������������������       ��2�s@:             X@������������������������       ���%�t_@`            @c@                           @`�5�#U�?P            �^@������������������������       ���	�H��?+            �P@������������������������       ����T�?%            �L@                           @�R �ΰ@�           �@                           �?{�HE	@k           ��@������������������������       ����0S�@�            �n@������������������������       �Bf�U	@�            �u@                           @�P
g(@l            @e@������������������������       ���*+A�?2            �Q@������������������������       �ܜ`�5d@:            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      s@     ��@     �@@      M@     �{@     �U@     $�@     �l@     H�@     �u@      7@      @     �h@     px@      *@      B@     �s@     @P@     ��@     �d@     `�@     @o@      .@      @     @a@     @g@      @      ;@     `i@     �H@     �o@      `@     �m@     `b@      *@             �^@      d@      @      :@      e@      @@     �m@     �Z@     `j@     �X@      (@              B@     �D@              @     �K@      @     �[@      "@     �V@      3@      @             �U@      ^@      @      5@     �\@      ;@     �_@     @X@     @^@     �S@      "@      @      0@      9@       @      �?      A@      1@      0@      7@      ;@     �H@      �?      @       @      4@              �?      4@      *@      &@      "@      ,@      ?@              �?      ,@      @       @              ,@      @      @      ,@      *@      2@      �?      �?     �M@     �i@      @      "@     �[@      0@      �@     �B@     �s@     �Y@       @              <@     �Y@      @      @      D@       @     v@      .@     `e@     �J@                      ,@      @@                      1@             �e@      @     �K@      &@                      ,@     �Q@      @      @      7@       @     `f@      &@      ]@      E@              �?      ?@     �Y@      @      @     �Q@      ,@     �c@      6@     `b@      I@       @      �?       @      3@                      (@      @     �F@      @      <@      ,@       @              7@      U@      @      @     �M@       @     �\@      2@     �]@      B@              (@     �Z@      a@      4@      6@     �`@      6@     �p@     �O@     �o@     �W@       @      @      :@      A@      @      @      =@      @     @]@      0@     �Y@      >@              @      5@      >@      @      @      6@      @     �P@      ,@      J@      :@              �?      ,@      &@      @              (@              A@      @      (@      @              @      @      3@              @      $@      @      @@      &@      D@      5@                      @      @                      @             �I@       @      I@      @                      @      �?                                      A@       @      8@      �?                      �?      @                      @              1@              :@      @               @     @T@     �Y@      0@      .@      Z@      2@     �b@     �G@     �b@      P@       @       @      R@     �V@      .@      &@     �V@      2@     �V@      E@     �Y@     �G@      @      @      ?@     �C@      $@      @      >@      @      >@      $@     �K@      7@      @      @     �D@      J@      @      @     �N@      ,@      N@      @@      H@      8@      @              "@      (@      �?      @      *@              N@      @      H@      1@      �?               @                              $@              >@              9@      @      �?              @      (@      �?      @      @              >@      @      7@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�{���N@�	           ��@       	                    �?���,@           ,�@                           �?��� �@1           �}@                            @�{�x�@y            @g@������������������������       ���9��@S             _@������������������������       �* eK�@&             O@                            �?J�
%�g@�            0r@������������������������       ��}��q@Z            �a@������������������������       ���y[i@^            �b@
                           �?��z�	�@�           p�@                           @���f@           @{@������������������������       ��ӊ���@l            �e@������������������������       ��\Dі @�            Pp@                          �7@��E �@�            �s@������������������������       �����[ @�            �o@������������������������       �_�J�y�@(            �N@                           �?p�9�8U@�           ��@                          �8@�/1�)
@�           ȑ@                          �4@T�4�a�	@�            �@������������������������       �X9Χ�e	@�            �x@������������������������       �Ǔ�x%	@�            `w@                           �?o?�w�/
@�             w@������������������������       ���Ӄ�@D            @X@������������������������       ���"��
@�            q@                          �2@��P�@�           0�@                           @̠ζ[@           |@������������������������       ����.6�@p             h@������������������������       �D����� @�             p@                           �?e��@�           ,�@������������������������       �nP]	@.            �Q@������������������������       �����S�@�           �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     ��@      =@      N@     Py@     �U@     ��@      k@     0�@      v@     �C@             @R@      h@      �?      $@     �X@       @     p}@      D@     `n@     �T@      @              E@     �X@      �?      @     �N@       @     @Y@      5@      W@     �H@      @              .@      >@                      7@              K@      @      G@      .@                      (@      1@                      4@              >@       @      =@      ,@                      @      *@                      @              8@      �?      1@      �?                      ;@      Q@      �?      @      C@       @     �G@      2@      G@      A@      @              ,@      A@      �?       @      ,@              3@      @      <@      4@      @              *@      A@              @      8@       @      <@      (@      2@      ,@                      ?@     �W@              @      C@      @      w@      3@     �b@      A@       @              ,@      P@              @      :@      @      l@      ,@     �Q@      .@                       @      8@               @      ,@      @     @T@      @      >@      "@                      @      D@               @      (@              b@      &@      D@      @                      1@      ?@                      (@       @      b@      @     @T@      3@       @              1@      ;@                      @             �_@       @      N@      (@       @                      @                      @       @      2@      @      5@      @              3@      l@     �w@      <@      I@      s@     �S@     ��@      f@     ��@     �p@     �@@      2@     @^@     �e@      4@      >@     �c@      J@      a@     @[@     �b@     �b@      :@      $@     @V@     @_@      @      ;@      [@      >@      Z@     �I@      ]@     �U@      0@      @     �F@      D@      @      $@     �K@      *@      S@      ?@     �N@      G@      @      @      F@     @U@              1@     �J@      1@      <@      4@     �K@      D@      $@       @      @@     �H@      ,@      @      H@      6@      @@      M@      @@      O@      $@       @      @      (@      �?              5@      @      "@      ,@      "@      4@       @      @      <@     �B@      *@      @      ;@      3@      7@      F@      7@      E@       @      �?     �Y@     �i@       @      4@     �b@      ;@     �|@     �P@     �w@     @^@      @              ,@     �N@               @      ;@      @     �h@       @     �Z@      >@                      @      @@              �?      &@      @     @V@      @      <@      .@                      @      =@              �?      0@              [@      �?     �S@      .@              �?     @V@      b@       @      2@     �^@      8@     0p@     �M@     @q@     �V@      @      �?      "@      (@               @      @      @      @      "@      &@      @                      T@     �`@       @      $@      ]@      4@     �o@      I@     �p@      V@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ\�qShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?T`-�@�	           ��@       	                    �?H�U�@           ��@                          �3@0B�d��@�            �@                          �1@Q���P@�            �q@������������������������       ���X,(�?Q             ^@������������������������       ��H/�J<@d            �d@                           �?~��fw@@�            �v@������������������������       ��/��J@_             b@������������������������       ��E����@�             k@
                           �?r��g@k           8�@                          �5@,�P,@�            �k@������������������������       ��@t@L            @]@������������������������       �7,3��@N             Z@                          �8@��ac4@�            �t@������������������������       �����f@�             q@������������������������       �z)A8;�?              M@                           @O�o,|@�           <�@                           �?+�3���	@�           T�@                           @]��ф�	@f           Ȃ@������������������������       �n���|@�            0q@������������������������       ����9j�	@�            `t@                           �?)hhd[	@�           ��@������������������������       ����@:            �X@������������������������       �����U'	@L           Ќ@                           @���;�@�           $�@                          �5@T@_��;@�           ��@������������������������       �Ʊ��ڸ@�           ȅ@������������������������       �zL�h�@�             w@                            �?�i�`Q	@             >@������������������������       ���1�@	             1@������������������������       �ZX�J��@
             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     �@      A@     @Q@     �{@     �X@     Ў@     `k@     ��@     �w@      =@      �?     �R@     `e@      �?      $@     �Y@      2@     pz@      F@     �p@     �S@      @      �?      C@      T@      �?      @      O@      &@      p@      >@     �\@     �D@                      $@     �A@                      0@      �?      a@      .@     �O@       @                      �?      (@                      @             �P@      @      8@      @                      "@      7@                      "@      �?     �Q@      "@     �C@      @              �?      <@     �F@      �?      @      G@      $@     �^@      .@      J@     �@@              �?      1@      6@      �?      @      2@      @      <@      &@      3@      4@                      &@      7@              @      <@      @     �W@      @     �@@      *@                     �B@     �V@              @     �D@      @     �d@      ,@      c@     �B@      @              5@      D@              @      ?@              E@      &@     �J@      2@       @              @      4@               @      $@              @@      @      B@      @                      ,@      4@              �?      5@              $@      @      1@      *@       @              0@     �I@                      $@      @     �^@      @      Y@      3@      �?              0@      F@                      $@              ]@      @     �P@      0@                              @                              @      @             �@@      @      �?      *@     �m@     `y@     �@@     �M@      u@      T@     ��@     �e@     P~@     �r@      :@      *@     �e@     p@      ;@     �E@      n@     �M@     @k@     �b@      l@     �h@      4@      @     �N@     @Z@      .@      ,@     �X@      9@      N@     �J@     @R@     �T@       @      @      <@     �H@      "@              J@      .@      :@      0@     �A@     �D@              �?     �@@      L@      @      ,@     �G@      $@      A@     �B@      C@      E@       @       @     �[@      c@      (@      =@     �a@      A@     �c@      X@     �b@     �\@      (@      �?      "@      @              &@      2@      @      $@      .@      ,@      *@      �?      @     �Y@     �b@      (@      2@      _@      ?@     �b@     @T@      a@     �Y@      &@             �P@     �b@      @      0@     @X@      5@     �u@      :@     Pp@     �Y@      @             @P@     `b@      @      (@     �V@      2@     Pu@      9@     0p@     �X@      @              7@     �X@       @      @      E@       @     `o@      ,@     @h@      J@      @              E@     �H@       @      @     �H@      $@     �V@      &@     @P@     �G@                       @       @       @      @      @      @      @      �?       @      @                                       @      @       @      @       @              �?      @                       @       @                      @               @      �?      �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ1 �hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Hٻ�wl@�	           ��@       	                   �3@0���H�@�           8�@                          �2@��I@�           ��@                           �?/���e@+           P}@������������������������       ��H��@g             e@������������������������       ���M+�@�            �r@                           �?�JsC�@�            �l@������������������������       �]��s �@_            �c@������������������������       �j��T7@.            �R@
                           �?N��l	@�           ��@                          �;@a)M�s�@           |@������������������������       ��- Ǒ@�            �u@������������������������       �i ��	@9             Z@                          �8@-͙7(�	@�           |�@������������������������       �L�$g�	@�           ؂@������������������������       �Z�ކU<
@)           @|@                           �?�Y���!@4           ��@                            �?���Y� @_           ��@                          �7@'�-@�            �q@������������������������       �a�Dj2 @�             m@������������������������       ��$��S@             �H@                            @X��;1�?�             p@������������������������       �.(l����?o            �e@������������������������       ��:_"�?:             U@                           @"�ycG@�           D�@                           @�<Qn!@           `�@������������������������       �����-@�             r@������������������������       �*Ǔ3��@\           P�@                            �?��U	g@�            Pt@������������������������       ���,�}f@*             S@������������������������       �����
@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Ps@     ��@      @@     �N@     �|@     @U@     ؏@      m@     ��@     �t@      A@      2@     �j@      t@      7@      G@     �t@      O@     �w@     `g@     �v@     `l@      >@       @     �F@      Y@      �?      "@     �U@      0@     `f@     �N@     �]@     �S@      @      �?     �@@     �P@              @      R@      @     ``@     �B@     �R@     �F@       @              @      2@                      8@              Q@       @      D@      &@              �?      <@      H@              @      H@      @     �O@     �A@      A@      A@       @      �?      (@      A@      �?      @      .@      *@      H@      8@      F@     �@@       @      �?      @      7@      �?      @      *@      *@      =@      ,@      5@      =@       @              @      &@              �?       @              3@      $@      7@      @              0@     �d@     �k@      6@     �B@     �n@      G@     `i@     �_@     �n@     �b@      :@       @     �G@     �R@      @       @     �N@      @     @W@      9@     �U@      B@      @             �A@      L@      @      @     �H@       @      V@      0@     @Q@      2@      @       @      (@      3@              @      (@      @      @      "@      1@      2@       @      ,@      ^@      b@      3@      =@      g@      D@     �[@     @Y@      d@     @\@      3@      @     �P@     �U@      (@      3@      `@      6@     �O@      C@     @Y@     �L@      @      $@      K@     �M@      @      $@     �L@      2@     �G@     �O@     �M@      L@      (@             @X@     �j@      "@      .@      `@      7@     �@      G@     �z@     �Z@      @              0@     @Q@                      <@      @     0p@      &@     �`@      .@                       @      E@                      7@      @     �]@      @      Q@      &@                      @     �@@                      3@      �?     @\@      �?      K@       @                      @      "@                      @      @      @      @      ,@      @                       @      ;@                      @             �a@      @     �P@      @                      @      :@                      @             @V@      @     �D@       @                       @      �?                      �?             �I@      �?      :@       @                     @T@     @b@      "@      .@     @Y@      0@     �w@     �A@     Pr@     �V@      @              I@     �\@      @      @      R@      "@     �r@      1@     �j@      N@      @              8@     �G@       @      �?      6@      "@     �V@      (@     �L@      7@      @              :@     �P@       @       @      I@             �i@      @     �c@     �B@                      ?@      @@      @      (@      =@      @     @T@      2@     �S@      ?@      �?              "@      @              @       @      �?      >@      @      4@       @                      6@      ;@      @      "@      ;@      @     �I@      ,@      M@      =@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ|�<%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�g�HR@�	           ��@       	                    �?발��@�           ��@                           �?E�z��1@�           ��@                            �?z��}�@~             j@������������������������       ��#m��@S            �`@������������������������       �~��-�/@+             S@                            �?��(WCx@:           P~@������������������������       ��2(H�@^            `b@������������������������       ����d�@�             u@
                          �5@-��l�>	@�           ��@                           �?$jg��1@�           ��@������������������������       �q��O�@J           0�@������������������������       ��W�K�?@�            �m@                           @�j�r޽	@           x�@������������������������       ���X	��	@�           ��@������������������������       ��G<D�p@P            �_@                          �4@i�M��@2           ��@                           �?߀�c*}@D           x�@                            �?pޣ��?�            �t@������������������������       ���"���?}            @g@������������������������       �_�N�y��?_            �b@                           @2+���@h            �@������������������������       �Y	���@a           ��@������������������������       ��r�u�@             ,@                          �<@Ć\fM@�           �@                            �?����B�@�            �@������������������������       ��/� @]            �b@������������������������       ��w����@U           H�@                            �?5+��q�@<            @X@������������������������       ���6���@            �F@������������������������       �"̳(�@             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     @r@     (�@      @@     �K@      @     �T@     `�@     �k@      �@     �t@     �@@      .@     `j@     �t@      8@      C@     �v@     �M@     `v@     �g@     Pz@     @l@      9@      �?      O@      [@       @       @     @V@      @     �c@      :@     `e@      N@      @      �?      4@      >@                      >@              N@       @     �I@      &@      @      �?      .@      0@                      (@              C@      �?     �A@      &@      @              @      ,@                      2@              6@      �?      0@                              E@     �S@       @       @     �M@      @     �X@      8@      ^@     �H@      �?               @      @@               @      @      �?      ;@      @     �K@      (@                      A@      G@       @      @      K@       @      R@      3@     @P@     �B@      �?      ,@     �b@     `l@      6@      >@     q@      L@     �h@     �d@     @o@     �d@      4@      @     �K@     @[@      $@      *@     `a@      &@     �`@     @R@     �^@      T@      @      @      G@     �R@      "@      "@     �\@       @     �P@     �H@     @S@      K@      @              "@      A@      �?      @      8@      @     �P@      8@      G@      :@              "@     �W@     �]@      (@      1@     �`@     �F@     @P@      W@     �_@     �U@      0@      @     @T@     �X@      &@      1@     @\@     �D@      M@     �O@     �[@      S@      (@      @      *@      3@      �?              5@      @      @      =@      0@      $@      @             @T@     �j@       @      1@     �`@      8@     0�@      =@     �y@      [@       @              A@     @Z@       @      @     �I@      @     �y@       @     �j@      G@                      $@      B@              �?      $@             �h@      @     @P@      (@                      @      1@                      "@             �Z@             �B@      &@                      @      3@              �?      �?              W@      @      <@      �?                      8@     @Q@       @      @     �D@      @     @j@      @     �b@      A@                      8@      Q@       @      �?     �D@      @     �i@      @     `b@      >@                              �?              @                      @              @      @                     �G@     @[@      @      (@     �T@      3@     �i@      5@     �h@      O@       @              B@     �X@      @      $@     �N@      1@     �h@      4@      f@     �E@       @               @      *@       @              &@      @     �K@       @      C@      2@                      <@     @U@      �?      $@      I@      *@      b@      2@     `a@      9@       @              &@      &@      @       @      6@       @      @      �?      3@      3@                       @      "@                      @       @      �?              $@      "@                      @       @      @       @      0@              @      �?      "@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?/7 t�0@�	           ��@       	                    �?3L<�C�@           L�@                            �?06M<mC@C           0�@                          �;@���@_            �c@������������������������       �,Xf��@V            �a@������������������������       �Q|���� @	             2@                            �?$���h@�            �v@������������������������       ���:���@W            �a@������������������������       �����s�@�            `k@
                          �5@���ix�@�           h�@                           �?B�r8� @J           H�@������������������������       �R��w� @�            @r@������������������������       ����TmB�?�            �l@                           �?D9,��@�            �h@������������������������       �@�^�q(@J            �Z@������������������������       �&;���2@;            @V@                           �?R��M�@�           �@                           @>�$/*	@�           t�@                           �?��77 �	@�            `m@������������������������       ��UtL�@!            �L@������������������������       �g�;.	@u            @f@                           �?ݼ�bx�@+           ��@������������������������       �\�Q�@�            �t@������������������������       �ڐڭhN	@c           H�@                           @�f�#b@�           d�@                           @:i��7
@�           `�@������������������������       �� O�[�@           py@������������������������       ��B6/��@�            Pq@                          �4@WS<�?�@           h�@������������������������       ����j}�@           P{@������������������������       ����:FN@           �{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pr@     �@      5@     �K@     `~@      Q@     �@     `i@     ��@     �y@     �@@      �?     @Q@     �c@      @      *@     �^@      "@     �|@      C@     �p@     �T@       @      �?      D@      U@      @      &@     @R@      @     �[@      <@     �[@      G@      @      �?      ,@      @@              @      4@       @      =@      @      F@      @      �?              "@      ;@              @      .@              =@      @      F@      @      �?      �?      @      @                      @       @                                                      :@      J@      @      @     �J@       @     �T@      8@     �P@     �C@      @              .@      ,@       @       @      2@              ;@      $@      =@      4@      @              &@      C@       @      @     �A@       @     �K@      ,@      C@      3@                      =@     @R@      �?       @     �H@      @      v@      $@     �c@     �B@      @              5@      M@               @     �B@       @     �q@      @     �W@      0@      @              $@     �B@               @      ;@       @     �c@      @      E@      &@                      &@      5@                      $@              _@       @     �J@      @      @               @      .@      �?              (@      @     �Q@      @     �N@      5@                      @      @                      @             �E@      �?      @@      .@                      @       @      �?              @      @      <@      @      =@      @              1@      l@     Px@      0@      E@     �v@     �M@     ��@     �d@     `~@     `t@      9@      0@     �^@     �f@      *@      2@     `g@      =@     @_@      W@     �b@     `d@      2@      @      =@      ?@      @      @     �@@      "@      0@      7@      H@      9@      @      �?      @      $@      @              1@                       @      @      (@      �?      @      9@      5@              @      0@      "@      0@      5@     �E@      *@      @      "@     �W@     �b@       @      .@     @c@      4@     @[@     @Q@     �Y@     @a@      (@              8@     �N@               @      N@       @      M@      3@     �B@     �L@      @      "@     �Q@     �V@       @      @     �W@      2@     �I@      I@     �P@     @T@      "@      �?     @Y@     �i@      @      8@      f@      >@     �{@     @R@     �t@     `d@      @      �?     �D@     �Y@              @     �X@      5@     �e@     �F@     �\@      S@      @              8@     �N@              @     �M@      .@     �T@      B@     �R@     �G@       @      �?      1@      E@              �?     �C@      @     �V@      "@     �D@      =@       @              N@      Z@      @      1@     �S@      "@     �p@      <@     �k@     �U@      @              5@     �E@       @      @      3@      �?     �d@       @      `@     �F@                     �C@     �N@      �?      ,@      N@       @     @Y@      4@     �V@      E@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @*kv�v@�	           ��@       	                    �?6��Ħ 	@o           :�@                           �?L�(l�f@�           `�@                          �8@B�"C@           �{@������������������������       �����@�            0t@������������������������       ��*-TL@L            �^@                          �3@f�}
�X@}            �i@������������������������       �?)�E@:             Y@������������������������       �\�w�,�@C            �Z@
                          �:@f��6H�	@�           D�@                           �?��QҘ	@           ��@������������������������       ���T�s	@           �{@������������������������       ��)mP�@�           h�@                            @�X(%
@�            �r@������������������������       ����a�	@v            @g@������������������������       ��4���?	@H            �[@                           @�5�#)@T           ��@                          �=@��Q )@�           ,�@                            @_Ae0��@�           ��@������������������������       �l@j`�@}           @�@������������������������       �G�(�~�?\            @c@                            �?#���Z@            �D@������������������������       ��#�A=)@
             1@������������������������       �����_/@             8@                            @��K��@e           �@                           @h�܎L-@            y@������������������������       ��.���@�            @r@������������������������       �"m����@L            �[@                           �?������@Z            �a@������������������������       �ɴ7mpT@.            �Q@������������������������       ��{�f�@,             R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     `�@     �B@     �M@     �{@     �T@     ��@     `j@     p�@     0x@     �@@      3@     @k@     �s@      6@     �E@     �r@      Q@     0w@     �e@     �w@     �p@      ?@              Q@     @U@      @       @      R@      "@     @e@      <@     �a@     �P@      @              K@     �Q@      @       @     �L@      @     @U@      8@      W@     �H@      @             �@@      H@      @              A@      @     @S@      2@     �R@      :@      @              5@      7@               @      7@               @      @      1@      7@                      ,@      ,@                      .@      @     @U@      @      I@      2@       @              (@      @                      @             �@@      �?      @@      (@                       @       @                      &@      @      J@      @      2@      @       @      3@     �b@      m@      3@     �D@     `l@     �M@      i@      b@     �m@     �h@      9@      @     �\@      i@      $@      A@     �f@     �E@     �f@      ]@     �j@     �`@      5@       @     �D@      V@      @      $@     �L@      (@     �L@     �K@      L@      J@      "@      @     @R@      \@      @      8@     �_@      ?@      _@     �N@     �c@     �T@      (@      *@      B@     �@@      "@      @      F@      0@      4@      =@      7@     �O@      @      $@      *@      3@      @      @     �@@      .@      $@      6@      *@     �D@       @      @      7@      ,@      @       @      &@      �?      $@      @      $@      6@       @             �S@     �m@      .@      0@      b@      ,@     �@      C@     0{@     �^@       @             �F@     �d@      @       @     �V@      @     �|@      9@     r@     �Q@      �?             �D@     �d@      @      @      S@      @     `|@      6@     �q@     �P@      �?              B@     �c@      @      @      P@      @     `x@      4@     �k@     @P@      �?              @      "@                      (@              P@       @      N@       @                      @                      @      ,@              @      @      "@      @                      �?                              @              @              @      @                      @                      @      $@              �?      @      @                             �@@     @R@      $@       @      K@      @     `b@      *@     @b@     �J@      �?              >@     �M@      @      @     �E@      @      X@      (@      \@      >@      �?              0@      H@      @      �?      <@      @     �S@      @     @V@      ,@      �?              ,@      &@              @      .@       @      2@      @      7@      0@                      @      ,@      @      �?      &@       @     �I@      �?      A@      7@                               @      �?      �?      @       @      >@              1@      @                      @      @       @              @              5@      �?      1@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�BChG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��sB�P@�	           ��@       	                    �?����J�@~           N�@                           �?�@��w@�           X�@                           �?����@~             i@������������������������       ����2��@8            �W@������������������������       ��bT3�}@F            �Z@                           �?]�)��@)           0|@������������������������       �����@�            �p@������������������������       �Nb]��@z            @g@
                           �?,h,��c	@�           p�@                           @�.-o�	@�           ��@������������������������       �����dz	@�           P�@������������������������       �Y%7=g@             ;@                            @Ψ O�@           �z@������������������������       ������~@�            Pr@������������������������       ��?b:@S             a@                          �7@�\�I@*           ��@                          �1@��
�@0           l�@                           @�O�!!; @�            pv@������������������������       �ƄI�� @�             r@������������������������       �����(�?*            �Q@                           �?vK�C�@W           ��@������������������������       ����w�p�?�            pr@������������������������       �)<��@�           h�@                          �<@4�^<�t@�            px@                            @%M�P��@�            �r@������������������������       ���֞�@�             n@������������������������       ��;����@%             N@                           @J�x�@8            �V@������������������������       �ـ�Xw@            �A@������������������������       �;��a��@#            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     ��@      @@      K@     P|@     �T@      �@     �j@     P�@     �u@      =@      4@     �i@     �u@      4@      E@     ps@     �Q@     �v@     `f@     �x@      n@      6@      �?     �Q@     �V@       @       @     @T@      @      d@      =@     �a@      N@      @      �?      7@      ;@                      8@              Q@      @      C@      ,@       @      �?      *@      "@                      ,@             �A@      �?      ,@      @                      $@      2@                      $@             �@@       @      8@      @       @             �G@     �O@       @       @     �L@      @      W@      :@     @Z@      G@      �?              ?@      G@       @       @      D@      @      @@      4@     �H@      A@                      0@      1@                      1@      �?      N@      @      L@      (@      �?      3@      a@     �o@      2@      A@     �l@     �P@     �i@     �b@     �o@     �f@      3@      3@     �Y@     �d@      ,@      8@     @f@     �J@     �`@     �[@      f@      b@      2@      (@      Y@     `d@      ,@      8@     �e@     �J@     �`@     �Z@     �e@     �a@      *@      @       @       @                      @                      @      @      �?      @             �A@     �V@      @      $@      J@      *@      R@      D@      S@      B@      �?              ?@     �H@      @      "@      F@      &@     �B@      ;@     �L@      8@      �?              @     �D@      �?      �?       @       @     �A@      *@      3@      (@              �?     �S@     �n@      (@      (@     �a@      *@     ��@      A@     �{@      [@      @              M@     �h@      "@      @     �W@      $@     �@      "@     u@     @P@      @              @      E@              @      7@             `f@       @     �V@      $@      @              @     �B@               @      6@             �`@             @S@      @      @                      @              �?      �?              G@       @      *@      @                     �I@     �c@      "@      @     �Q@      $@      u@      @     �n@     �K@      @              $@      F@      �?              *@      �?     �b@      �?     �Q@      @                     �D@      \@       @      @      M@      "@     �g@      @      f@     �H@      @      �?      5@     �H@      @      @      H@      @     @T@      9@     �[@     �E@      �?      �?      ,@      B@      �?      @      >@      @      R@      8@     @V@      :@      �?      �?      (@      A@              @      8@      @      D@      4@      T@      7@      �?               @       @      �?      �?      @              @@      @      "@      @                      @      *@       @       @      2@              "@      �?      5@      1@                      �?      @       @       @      @              @      �?      $@      @                      @       @                      .@              @              &@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Y4�w@�	           ��@       	                   �;@�����@�           ��@                           �?����@�           ��@                           �?��{ar	@S           �@������������������������       ��]�0v�@G           p@������������������������       �+��|��	@           �@                           �?�A!$��@i           8�@������������������������       ��P�G�	@j             d@������������������������       �tnE���@�            `x@
                           �?(3�B�	@�            �v@                            �?�"i�8@8            @W@������������������������       ����h@"             K@������������������������       ���Mc��@            �C@                            @8��V[
@�            �p@������������������������       �}&dF��	@U             c@������������������������       ����U�g	@D             ]@                          �7@��	�	@           ��@                           �?x�8Rj�@           �@                           @�:�1:2 @           {@������������������������       �s��`�?�            0q@������������������������       ���~\F�@^            �c@                          �1@B_+��@           @�@������������������������       ��S��:s�?r            �g@������������������������       �S��p@�           `�@                           @Ù:l5I@�            `x@                           @#�
NQ@�            �l@������������������������       �qvq�2�@H             ^@������������������������       ����:�@H            �[@                           �?�ޯ%@�@i             d@������������������������       ������@/            �R@������������������������       ���6v@:            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      t@     0�@      ?@     �N@     p|@     @U@     ��@     �k@     ��@     �t@     �B@      1@     �m@     Pt@      :@     �H@     �s@     @P@     �v@     �f@     �y@     �l@      >@      "@      h@     @q@      1@      C@     q@     �F@     pt@     �b@     �v@     `e@      >@      "@      b@     �h@      .@      >@      j@      A@     @g@     �[@      o@     @_@      =@              A@      U@      �?      ,@     �T@      @      V@     �A@     @Y@      H@      "@      "@     �[@     �\@      ,@      0@     �_@      <@     �X@     �R@     `b@     @S@      4@             �G@     �S@       @       @      P@      &@     �a@      C@     �\@      G@      �?              $@      *@              �?      (@       @     �Q@      �?     �E@      "@                     �B@     @P@       @      @      J@      "@     �Q@     �B@      R@     �B@      �?       @      G@     �H@      "@      &@      F@      4@      A@      A@      H@      M@                      @      &@       @      @      0@       @      &@      "@      .@      2@                       @       @                      $@       @      @      "@      $@      "@                      @      @       @      @      @              @              @      "@               @      D@      C@      @       @      <@      2@      7@      9@     �@@      D@              @      4@      (@       @      @      2@      &@      "@      0@      :@      <@              @      4@      :@      @      @      $@      @      ,@      "@      @      (@              �?      U@      l@      @      (@     @a@      4@     h�@     �C@     `y@     @Z@      @             �N@     �e@      @      "@      W@      (@     ��@      0@      s@     �O@      @              (@     �H@              �?      :@      @     �l@      @      X@      (@      @              @      8@                      (@      @     @d@       @     �O@      @                       @      9@              �?      ,@             �P@      �?     �@@      @      @             �H@      _@      @       @     �P@      "@     �r@      *@     @j@     �I@      @                      4@               @      (@              V@      �?     �M@      @                     �H@      Z@      @      @      K@      "@     �j@      (@     �b@     �F@      @      �?      7@      J@      �?      @      G@       @     �V@      7@      Y@      E@              �?      (@      B@              �?      8@      �?      Q@      @      O@      4@              �?       @      2@              �?      &@      �?     �I@      �?      ?@      @                      $@      2@                      *@              1@      @      ?@      1@                      &@      0@      �?       @      6@      @      7@      2@      C@      6@                      @      (@              �?      @      @      *@      @      4@      @                      @      @      �?      �?      .@      @      $@      &@      2@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJGo#5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �1@ޔ��Ia@�	           ��@                          �0@_,yϦS@�           0�@                           @_T��4@            �j@                           �?�F�D�@d            @e@������������������������       �Ĉp�I@6            �Y@������������������������       �U��FV@.            �P@������������������������       ��&��1��?            �F@                            @���!@           �x@	       
                    �?��G��g@�            �q@������������������������       �3.EF� @Z            �a@������������������������       ��30	G @b            @b@                           �?���G@F            @\@������������������������       �n�&�(@            �I@������������������������       �U�Z���@*             O@                           @@�!���@-           Ʃ@                          �;@J��U�@	@�           �@                          �4@8beᏼ@           ̙@������������������������       ���^�@�           ��@������������������������       �z�r��@s            �@                           �?b��	�I
@�            �t@������������������������       �_��*��@;            @W@������������������������       �{�-d[�
@�             n@                          �8@ ���@Z           ��@                           �?�O;��0@�           `�@������������������������       ��e�@T           �@������������������������       ��;.�@?           �~@                          �<@��:Q�@�            `s@������������������������       ���Cq�@�            `j@������������������������       ��)�R@@            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     �q@     ؁@      @@     �M@     �z@     �Q@     ��@     @o@      �@     �v@      C@              ,@     �T@      �?      @     �H@      �?     0q@      <@     ``@      <@                      @     �C@              �?      8@             �V@      @      D@      (@                      @      8@              �?      8@              Q@      @      B@      $@                       @       @                      ,@             �F@       @      :@      @                      �?      0@              �?      $@              7@       @      $@      @                              .@                                      6@       @      @       @                      &@     �E@      �?      @      9@      �?      g@      6@     �V@      0@                      @      =@              @      2@      �?     `a@      &@     �P@      &@                      @      ,@              @      (@      �?      Q@      @      <@      @                      @      .@                      @             �Q@      @     �C@      @                      @      ,@      �?              @              G@      &@      8@      @                       @      "@      �?              �?              9@      "@      �?      @                      @      @                      @              5@       @      7@       @              1@     �p@     �~@      ?@      K@     �w@     @Q@     `�@     �k@     �@     0u@      C@      1@     �h@     Pr@      7@      E@     �p@      M@     �s@      g@     �s@     �m@     �@@      "@     �c@     @o@      ,@      <@     `m@     �F@     r@     �b@     �q@     �d@      9@      @     �D@     �Q@       @      @     �R@      ,@      a@     �O@      `@      R@      &@       @     @]@     �f@      (@      5@      d@      ?@      c@     �U@     @c@     �W@      ,@       @     �D@     �E@      "@      ,@      B@      *@      :@     �A@      >@     �Q@       @      @      @      .@              @      @              @      (@      @      =@      @      @      A@      <@      "@      "@      >@      *@      3@      7@      9@      E@      @             �Q@     �h@       @      (@     �[@      &@     {@      C@     �t@     @Y@      @              I@     �d@      @       @     �T@      $@     pv@      2@     @m@     �P@      @              ;@     @T@       @      @     �K@      @     �d@      &@     �]@      F@      @              7@      U@      @       @      <@      @     `h@      @      ]@      7@       @              5@      ?@      @      @      ;@      �?     �R@      4@     �W@      A@                      $@      6@       @       @      $@      �?      L@      2@      R@      2@                      &@      "@      �?       @      1@              2@       @      7@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���X�R@�	           ��@       	                    �?*�*#jW@           ��@                          �<@��@9           �~@                          �:@Ǟ���@            z@������������������������       �7nq,�@�            �x@������������������������       ����}��@             :@                          @@@(�yl5�@*            �Q@������������������������       �k���@#             M@������������������������       �B�ޑL��?             *@
                          �8@�����@�           ��@                           �?�tB�Ǡ @�           ��@������������������������       ��s�� @�            @u@������������������������       ��i��%) @�            �p@                            @�M� �e@N             ^@������������������������       �*�|_e�@=             W@������������������������       ��E���?             <@                           @�DOZ#8@�           �@                          �6@�y5�	@X           ��@                           @��.O��@�           �@������������������������       �䷲^G@�           0�@������������������������       �X�ʢ6�@�           ��@                            �?1W��F	@           ��@������������������������       ����.B	@E           P�@������������������������       �����=�@:           ��@                           !@9r�8z�
@1            �R@                           �?l���	@#             J@������������������������       ����� �@             (@������������������������       ������V@             D@                           8@y;��@             6@������������������������       ��7���� @             &@������������������������       ��tc��@             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     @r@     ؁@      9@      G@     �}@     @W@     �@     @k@     P�@     0w@      ?@              R@     �f@       @      ,@     @W@      ,@     p{@      D@     Pq@      U@                      G@     @T@       @      &@      N@       @      \@      ;@     �X@     �H@                     �C@      Q@       @      @     �I@       @     @[@      :@     �W@      7@                      B@     �P@       @      @     �G@             �X@      8@     �V@      7@                      @      �?                      @       @      $@       @      @                              @      *@              @      "@              @      �?      @      :@                      @      (@              �?      @              @      �?      @      :@                              �?              @      @                              �?                              :@     �X@              @     �@@      (@     pt@      *@     @f@     �A@                      :@     �U@              @      9@      @     @r@      @      b@      7@                      "@     �J@              @      1@      @     �d@       @     �R@      (@                      1@     �@@                       @             @_@      �?     �Q@      &@                              *@                       @      "@     �A@      $@     �@@      (@                              *@                      @      "@      7@      "@      9@      $@                                                      @              (@      �?       @       @              2@     �k@     px@      7@      @@     �w@     �S@     X�@     @f@     P@     �q@      ?@      0@     �i@     x@      6@      >@     pw@     �Q@     �@     �d@      @     �q@      :@      $@     @X@     �m@      @      2@     @j@      :@     �y@     �T@     pr@     @a@       @      $@      P@      a@      @      &@     �a@      3@     `b@      R@     �[@     �U@      @             �@@     �X@       @      @     �Q@      @     �p@      $@      g@      J@      @      @     �[@     �b@      0@      (@     �d@     �F@     �`@     @U@      i@      b@      2@       @      N@     �R@      @       @     �R@     �A@     �M@      F@     �\@     �P@       @      @      I@     �R@      "@      @     �V@      $@     �R@     �D@     �U@     �S@      $@       @      *@      @      �?       @       @       @      "@      &@      @      @      @       @      "@      @      �?       @      @              "@      "@      @      �?      @      �?              �?               @      �?              @               @              �?      �?      "@      @      �?              @              @      "@       @      �?       @              @      �?                      �?       @               @      �?      @       @              @                                      @                      �?      �?       @              �?      �?                      �?      @               @               @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJhL^hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��շ<@�	           ��@       	                   �8@��6@           ��@                            �?7�^�g�@x           ��@                           @���w�@R           0�@������������������������       �j>c��f@�            pq@������������������������       ��}a��?�            �p@                           �?�8��!@&           �|@������������������������       �(Tv�Q�@�            `n@������������������������       ��-����@�            �j@
                          �<@#��@�             n@                           @���E�@^            �c@������������������������       �����Z@:            @X@������������������������       ��%Y"@$            �M@                           @����@6             U@������������������������       �W���_�@&             M@������������������������       �n�4�@             :@                          �2@��� T2@�           Ҥ@                           @�G���@�           ��@                           �?�5H��@�            �x@������������������������       �k�5f�`@�            `j@������������������������       �:l~�{l@p             g@                          �1@սr�lM@�            `p@������������������������       �!�o��?b            �b@������������������������       ��$�I&@A             \@                           @�Ӯ}��@�           \�@                          �:@�v�v�	@�           ��@������������������������       ����� N	@6           ��@������������������������       �ҝt�$
@�            �s@                           @Do/��*@�           P�@������������������������       ����� @_            �c@������������������������       ���F8@�           p�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@      �@      =@     �P@     `{@     @S@     0�@     @l@     �@     �v@      8@             @S@     �d@      @      "@      Y@      (@     �~@      F@      p@     �T@      @              K@     @_@      @      @     @Q@      @     �{@      @@     �j@     �I@      @              ?@     �O@      @      @      F@       @     @o@      (@     @]@      7@       @              >@      ;@       @      �?      9@       @      Y@      "@     @Q@      (@       @              �?      B@      �?       @      3@             �b@      @      H@      &@                      7@      O@               @      9@      @     �h@      4@     @X@      <@      �?              $@      ?@               @      3@      @      [@      @      I@      ,@                      *@      ?@                      @              V@      .@     �G@      ,@      �?              7@     �C@              @      ?@      @      H@      (@      E@      @@      @              1@      <@              �?      1@      @      B@      @     �@@      &@       @              1@      3@              �?      *@      �?      .@      @      .@       @       @                      "@                      @      @      5@      �?      2@      @                      @      &@              @      ,@       @      (@      @      "@      5@      �?              @       @              @      &@               @      @      @      0@      �?                      @                      @       @      $@              @      @              4@     �i@      x@      :@     �L@      u@     @P@     ��@     �f@     �@     �q@      2@      �?      A@      W@      "@      @     @P@       @     �h@      B@     @c@     �O@      �?      �?      >@     @P@       @       @     �D@       @     @Z@      A@     �O@      I@      �?      �?      4@     �A@       @      �?      ?@              B@      7@      @@      =@      �?              $@      >@              �?      $@       @     @Q@      &@      ?@      5@                      @      ;@      @      @      8@             �V@       @     �V@      *@                              0@               @      *@              P@      �?      I@      @                      @      &@      @      �?      &@              ;@      �?     �D@      "@              3@     `e@     @r@      1@      J@     q@     �O@     �u@     @b@     �x@     `k@      1@      2@     @]@      f@      *@      C@     �e@      I@     @b@     �^@     @f@      c@      *@      "@     @W@     �a@      @      ;@      `@      @@     @\@     �V@      b@      V@      "@      "@      8@      B@      @      &@      F@      2@     �@@      @@      A@      P@      @      �?      K@     �\@      @      ,@      Y@      *@      i@      8@     �j@     �P@      @      �?      @      6@       @      &@      9@      @      9@      (@      B@      (@                      H@     @W@       @      @     �R@      "@     �e@      (@     @f@     �K@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��� hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @C��<@�	           ��@       	                    �?"��ٻ@]           b�@                           �?�S|��	@�           x�@                           �?@P�k@y           ؂@������������������������       �V�i��@�            �i@������������������������       �}�I^�@�            �x@                           �?ciTo�	@i           �@������������������������       �{K���@�            Pt@������������������������       �6���
@�           ��@
                           �?s��"@{           ��@                          �<@L��*�@q             e@������������������������       �V�X�r8@j            �c@������������������������       ���!zȓ@             "@                          �4@���Ԩ@
           �z@������������������������       ��w� 
�@x            �h@������������������������       �oYF3@�            �l@                           @ӎ�� �@3           `�@                          �2@���@�           ܑ@                            �?}scC/�?           `x@������������������������       �P�^��?>            �Y@������������������������       ��6|� @�             r@                          �7@���d��@�           ��@������������������������       ��`=�
{@Z           ��@������������������������       ��Fp;�@�            �k@                           �?p0��4�@H           �@                          �6@��7^,�@�            �p@������������������������       �=Z��@m            �e@������������������������       ����V��@5            �W@                           @w����@�            0q@������������������������       �մ��@�             o@������������������������       �猵r;@             ;@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     p@     (�@      1@     �N@     0|@      V@     ��@     �l@     ؈@     �v@      =@      6@     `g@     `v@      $@      H@     `t@     �P@     `w@      g@     �v@     Pp@      7@      6@      b@     �p@      "@     �@@     �m@      M@      n@     @a@     �n@     @k@      4@      @      >@     @Y@              &@      X@      $@     �]@      D@     �[@     �S@      @      @      *@      =@                      ;@              J@       @     �J@      8@      �?      �?      1@      R@              &@     @Q@      $@     �P@      C@     �L@      K@      @      1@     �\@     `d@      "@      6@     �a@      H@     �^@     �X@     �`@     �a@      0@              A@     @P@               @      B@      @     �L@      6@      H@      G@      @      1@      T@     �X@      "@      ,@     �Z@     �E@     �P@      S@     �U@     �W@      (@             �E@     �W@      �?      .@     �U@      "@     �`@     �G@      ^@     �E@      @              &@      0@               @      *@      �?     �N@      @      I@      "@       @              &@      .@               @      *@      �?     �N@              H@       @                              �?                                              @       @      �?       @              @@     �S@      �?      *@     �R@       @      R@      F@     �Q@      A@      �?              @     �D@      �?      @      >@      �?      H@      3@      A@      .@                      =@     �B@              "@      F@      @      8@      9@      B@      3@      �?             �Q@     �k@      @      *@     @_@      5@      �@      G@     �z@     �Z@      @              D@      d@      �?      �?     �R@      $@     �|@      8@     �r@     �P@      @              @     �J@                      (@              i@      @     �X@      0@                              $@                       @             �Q@              0@      @                      @     �E@                      $@             ``@      @     �T@      (@                     �@@      [@      �?      �?     �O@      $@      p@      5@     �i@      I@      @              7@     �T@      �?      �?      B@      "@     @i@      *@     �`@      >@       @              $@      9@                      ;@      �?      L@       @     @R@      4@      �?              >@      O@      @      (@      I@      &@     �f@      6@      `@      D@      @              ,@      A@      @      "@      6@      @     �X@       @      K@      4@                      @      3@      @       @      ,@      �?     �R@       @      A@      ,@                       @      .@              �?       @      @      9@      @      4@      @                      0@      <@      @      @      <@      @     �T@      ,@     �R@      4@      @              ,@      8@      �?      @      :@      @     @T@      ,@      P@      1@                       @      @       @               @              �?              $@      @      @�t�bub�     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��&hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�Bx         
                   �1@�
?��d@�	           ��@       	                    @�X�jj�@|           P�@                            @ǒ46�?@m           ��@                           @����@           �x@������������������������       ��K$B�'@�             k@������������������������       ����Myi@y            `f@                           @z&��@k            �e@������������������������       �d��Ĵ@F            �[@������������������������       ��m=
��?%            �N@������������������������       �����z�@             3@                           �?�j�@+           ��@                           �?��K�*O@p           ��@                          �6@�W:�6%@           z@������������������������       �����YX@|            `i@������������������������       ��̸
�@�            �j@                            �?~�E��@o           ��@������������������������       �SFI/�x @X            �a@������������������������       � ���9@           �z@                           @�����@�           R�@                           �?
$&k m@           .�@������������������������       ��u��i�@m             h@������������������������       �Z�-.]^@�           \�@                          �3@+�`�(	@�             q@������������������������       �╌l��@$            �K@������������������������       ����?x	@�            `k@�t�bh�h5h8K ��h:��R�(KKKK��h��B`	        ,@     �q@     (�@     �B@     �L@     �z@     �X@     x�@     @k@     ��@     �v@      ?@      �?      .@     @S@              @     �I@      �?     �o@      6@     �`@      ;@      �?      �?      ,@     @S@              @     �H@             �n@      6@     ``@      7@      �?      �?      @     �M@              �?      C@             �e@      @     �V@      0@      �?              @      9@              �?      5@              [@      @      E@       @      �?      �?       @      A@                      1@             �P@      �?     �H@       @                       @      2@               @      &@             �Q@      .@      D@      @                      @      .@               @      $@             �@@      .@      ;@      @                      @      @                      �?              C@              *@       @                      �?                       @       @      �?      @               @      @              *@     �p@     �}@     �B@      J@     �w@     �X@     ��@     �h@     x�@     u@      >@             �R@     �`@      �?      "@      V@      ,@     Ps@      B@     �m@     @R@      @             �E@     �M@      �?       @     �M@      @     �S@      4@     �V@      I@      @              2@      ?@              @      .@       @      K@      @     �J@      4@                      9@      <@      �?      @      F@      �?      9@      *@      C@      >@      @              @@     @R@              �?      =@      &@     �l@      0@     �b@      7@       @              @      9@                       @      @     �P@              A@      @       @              =@      H@              �?      ;@      @     �d@      0@     �\@      2@              *@     �h@     @u@      B@     �E@     @r@      U@     �y@      d@      ~@     �p@      8@      @      f@     �q@      B@     �D@     �p@     @R@     @w@     �_@     �{@      m@      (@      @      8@      @@               @      A@      "@      ,@      &@     �F@      1@      �?      @      c@     �o@      B@     �C@     �l@      P@     `v@      ]@     �x@      k@      &@      @      3@      L@               @      ;@      &@     �D@     �@@      B@      ?@      (@              @      &@                      @      �?      *@       @      .@      @              @      0@     �F@               @      7@      $@      <@      ?@      5@      9@      (@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�#ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�Uߋ�M@�	           ��@       	                    �?z���V	@           p�@                          �:@�ϥ@+9@�           ��@                           �?��Mq�@C           p�@������������������������       �SB����@~            �i@������������������������       ����P�V@�             t@                           �?m)��@D            �[@������������������������       ���i��@            �B@������������������������       �y��>��@.            @R@
                           �?*��,)�	@z            �@                           �?�2�@�            pr@������������������������       ���D@Z            �a@������������������������       �5h����@c             c@                          �>@zS��
@�           ȅ@������������������������       ���3�	@�           ؃@������������������������       �m��@!             O@                           �?�?�S��@�           ڡ@                           �?�C65�@�           ȑ@                           @��SV�w @           pz@������������������������       ��	eH% @�            @p@������������������������       � ����M @m            `d@                            �?{2|�@�           X�@������������������������       �,�)u�z@c            �d@������������������������       �ɂ0y��@d           (�@                           �?4�ѱm@�           �@                          �9@�y<~�� @�            Pt@������������������������       �����
�?�            @q@������������������������       ��Ű�e3@            �H@                          �5@�?�%�@           ��@������������������������       ���d��Q@)           �}@������������������������       ���ٿnh@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@      r@     8�@      A@     �J@     `w@      V@     ,�@      m@     ��@     �w@      @@      4@     �c@     `n@      :@      @@     @m@     �H@     �l@     `a@     @p@     �j@      5@      @     �I@     �Y@      @      $@      S@      *@      _@     �F@     �]@     �S@      @      @      C@     �V@      @      "@      N@      $@      \@     �B@     �Z@     �J@      @      @      .@     �C@       @      �?      D@      @      I@      &@      <@      $@       @              7@     �I@      �?       @      4@      @      O@      :@     �S@     �E@      @      @      *@      *@       @      �?      0@      @      (@       @      *@      9@              @      &@      @                      @              @      @      �?      @                       @      @       @      �?      (@      @      @      @      (@      6@              *@     �Z@     �a@      5@      6@     �c@      B@     �Z@     �W@     �a@      a@      0@              5@      K@      @       @     �B@      @     �L@      2@     �J@      C@      @              @      >@      @      @      .@      @      ?@      "@      2@      4@      �?              ,@      8@               @      6@              :@      "@     �A@      2@       @      *@     �U@     �U@      2@      ,@     @^@     �@@      I@      S@      V@     �X@      *@      "@     �T@      Q@      .@      &@     @]@      @@      I@      P@     �U@     �U@      (@      @      @      2@      @      @      @      �?              (@      �?      (@      �?      �?     �`@     @s@       @      5@     �a@     �C@      �@     �W@     ��@     `d@      &@      �?      Q@      d@      @      (@     �T@      0@     z@     �A@     `n@     @V@      $@              ,@      I@               @      (@      @     �k@      @      V@      7@                      *@      ;@                      @      @      b@      @     �F@      0@                      �?      7@               @      @      �?     �S@      @     �E@      @              �?      K@     �[@      @      $@     �Q@      &@     @h@      =@     `c@     �P@      $@              .@     �C@                      2@             �A@      $@     �B@      "@      @      �?     �C@      R@      @      $@      J@      &@     �c@      3@     �]@     �L@      @              P@     `b@      @      "@      M@      7@     0x@     �M@     t@     �R@      �?              .@     �B@                       @      �?     �`@      @     �\@      $@      �?              .@      A@                      @             �_@      @     �U@      @                              @                      @      �?      @      @      ;@      @      �?             �H@     �[@      @      "@      I@      6@     �o@      J@     �i@      P@                      0@     �N@      �?      @      .@       @     @f@      6@      a@      >@                     �@@     �H@      @       @     �A@      ,@     @S@      >@     �Q@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��qWhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @o	r�8@�	           ��@       	                    �?�JU��@�           \�@                          �<@��`@�           �@                            �?%s�@�           �@������������������������       ��W#�@x             f@������������������������       �N����@           0{@                          �>@�5�V�6@#             O@������������������������       �NTu�@             E@������������������������       ��@p=�i@             4@
                          �1@�	2�z	@�           4�@                           �?����@i            �e@������������������������       �kB��B@*            �R@������������������������       �m���@?             Y@                            �?�Y��	@s           x�@������������������������       �ܦ�-�	@           py@������������������������       �qf'��	@q           8�@                           �?�d}��@5           l�@                            @�S��� @g           ȁ@                          �4@]���<@'           P}@������������������������       �y�N��?�            �r@������������������������       ��}B�`@i            �e@                           �?�
]	��?@             Y@������������������������       ��f�j�?%             N@������������������������       ��H7`~��?             D@                          �7@��v��A@�           ��@                           @�"�n�@@           ��@������������������������       �ۡխ@�           ��@������������������������       �1�D�/@�            `k@                           @�-��@�            �r@������������������������       �"�V<�A@w            �g@������������������������       �xB��@J            �\@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     Pr@     �@      6@      N@     �~@      P@      �@     @l@     0�@     `v@      >@      8@     �j@     �r@      ,@      G@     Pt@      G@     �w@      h@     �y@     `n@      :@              N@     �T@              @     �T@      @     �e@      8@     @f@      N@      @              K@      S@              @     �Q@      @     �e@      3@      e@      D@       @              2@      6@               @      ,@      �?      F@      @     �O@      @      �?              B@      K@               @     �L@       @      `@      ,@     �Z@      A@      �?              @      @              �?      (@              �?      @      "@      4@      �?               @      @              �?      @                      �?      "@      1@      �?              @      �?                      @              �?      @              @              8@     `c@      k@      ,@     �D@     @n@     �E@     �i@      e@     @m@     �f@      7@              0@      <@                      .@             �A@      7@     �E@      .@                      @      ,@                      @              4@      *@      $@      @                      &@      ,@                      "@              .@      $@     �@@       @              8@     `a@     �g@      ,@     �D@     `l@     �E@     `e@      b@     �g@      e@      7@       @      J@     �D@              *@      S@      ,@      I@     �M@     �F@     �F@      $@      6@     �U@     `b@      ,@      <@     �b@      =@     @^@     �U@     @b@     �^@      *@      �?     �S@     �j@       @      ,@     `d@      2@     @�@      A@     �z@     �\@      @              ,@     �Q@               @      @@       @     0q@      "@     �a@      5@       @              (@     @P@                      <@       @      k@      "@     �\@      4@       @              $@      B@                      $@             `d@      @      P@       @       @               @      =@                      2@       @      K@      @      I@      (@                       @      @               @      @              M@              <@      �?                       @       @               @      @             �B@              *@      �?                              @                      �?              5@              .@                      �?      P@      b@       @      (@     ``@      0@     Pu@      9@     �q@     �W@       @             �C@     �\@      @       @     @T@      ,@     �q@      (@     @j@     �I@       @              >@     �S@      �?      �?      F@      @     �l@      "@      d@     �B@       @              "@      B@      @      @     �B@      @      K@      @     �H@      ,@              �?      9@      >@      @      @      I@       @     �L@      *@     �R@     �E@              �?      .@      5@              @      ?@              G@      @     �H@      3@                      $@      "@      @              3@       @      &@      $@      9@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJE�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�� �@�	           ��@       	                    �?��Oس@           �@                            �?��s5f1@=           8�@                           �?�j���@^             a@������������������������       ��˪C:+@)            �N@������������������������       ���zo �@5             S@                           �?Lpk��@�            �w@������������������������       ������R@Y            �b@������������������������       �s�6���@�            @m@
                          �4@����@�           ؅@                           �?�55�r� @           �z@������������������������       ���Vʹ�@�            �m@������������������������       �
�ÈL�?}            �g@                          �=@�wm��#@�            �p@������������������������       �e�]PF@�             o@������������������������       ��׋�@             7@                          �4@u�ʱP@�           �@                            @k�r={@�           ��@                           @4M���@&           Ȋ@������������������������       ����@�            �v@������������������������       ���E��o@6           �~@                          �3@)n-�4@�            pt@������������������������       ��o>�dW@�            �o@������������������������       ���&?�@.            �R@                           @/�j�;	@�           ��@                          �9@ۍ4Ŕ�	@Z           ��@������������������������       �ٙuwK	@x           ��@������������������������       �ӕ�A5�	@�            �v@                           @�A���@g           @�@������������������������       �.��ۀ@Y           ��@������������������������       ��� ��@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     pq@     �@      ?@     �I@     �|@      U@     ��@     �n@     ��@      y@      ?@       @     @S@      c@      @       @     @]@      0@     �y@     �G@     �q@     �W@      @       @     �I@     �S@      @      @     �T@      �?     @X@      B@     �Z@      I@      @       @      "@     �@@              @      3@      �?      5@      @      B@      "@      �?       @      @       @                      (@              (@              4@      @      �?              @      9@              @      @      �?      "@      @      0@      @                      E@      G@      @      @      P@              S@     �@@     �Q@     �D@       @              .@      0@                      4@             �F@      @      B@      $@                      ;@      >@      @      @      F@              ?@      ;@     �A@      ?@       @              :@     @R@               @      A@      .@     �s@      &@      f@     �F@                      3@     �A@               @      0@              j@      @     @\@      ;@                      (@      6@               @      (@              ]@      @      H@      4@                      @      *@                      @             @W@             @P@      @                      @      C@                      2@      .@      [@      @     �O@      2@                      @     �B@                      0@      $@     @Z@      �?     �M@      ,@                      �?      �?                       @      @      @      @      @      @              5@     @i@     �x@      ;@     �E@     �u@      Q@     ��@     �h@     `@     s@      <@      @      N@     �e@      "@      *@     �]@      2@     pu@      Q@      o@     �]@      "@      �?      D@     @^@      @       @     @T@      $@     �p@     �I@      h@      S@      @      �?      9@     �M@      @      @      I@      @     �P@     �E@      Q@      B@      @              .@      O@              @      ?@      @     `i@       @     @_@      D@               @      4@      K@      @      @      C@       @     �R@      1@      L@      E@      @       @      2@      G@      @      @      9@      @      N@      (@     �E@     �A@                       @       @       @      �?      *@      @      ,@      @      *@      @      @      2@     �a@     @k@      2@      >@      l@      I@     �k@     @`@     �o@     `g@      3@      1@     �Y@      b@      ,@      7@     �c@     �D@      U@     �X@      `@     �`@      0@      "@     @Q@     �Y@      @      1@     �\@      5@     �J@      I@     �U@      M@      "@       @     �@@      E@       @      @     �D@      4@      ?@      H@      E@      S@      @      �?      D@     @R@      @      @     @Q@      "@      a@      @@      _@     �J@      @      �?      @@      R@      @      @     �P@      @      a@      >@      _@     �J@      @               @      �?      �?              @      @      �?       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ6�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�7=A�r@�	           ��@       	                     �?'�i1�@�           $�@                           �?�QH`@�            ps@                          �;@��WD%o@X            ``@������������������������       ���Tɯ�@P            �^@������������������������       �hJN�@             "@                           �?q�|��f�?s            �f@������������������������       �vP���?=             W@������������������������       ��� @6             V@
                            @�t"7��@*           ��@                            �?�ȿZk@`           ��@������������������������       ��H��@�            �w@������������������������       ����:�@�             k@                           @Ш؀s@�             t@������������������������       ��ݪ���@�            �l@������������������������       �˶�ؔG�?<            �V@                          �1@���?a@�            �@                           �?n`��?^@�            �v@                            @,>!�G)	@?            @X@������������������������       ����j_@"            �H@������������������������       ���9�@             H@                           @"��ـX@�            �p@������������������������       ���0�� @�            �j@������������������������       �^�\�V@             J@                           @�<����@�           *�@                          �:@�l-���	@u           ��@������������������������       ��"�-yY	@�           �@������������������������       ��n��	@�            �r@                          �7@�ڶ�9@K           `�@������������������������       ���НJ�@�           x�@������������������������       ��ǟT��@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     @s@     ��@      ?@      K@     {@     �T@     �@     @m@     ؇@     `v@      A@              W@     �e@      @      @     @V@      $@     �{@     �H@     �p@      V@       @              (@      I@       @              7@      @     �^@      "@     @R@      ,@      �?              (@      ;@                      .@       @      4@       @      C@      "@                      $@      :@                      ,@              4@       @     �B@      @                       @      �?                      �?       @                      �?       @                              7@       @               @      @     �Y@      �?     �A@      @      �?                      @                      @      �?      M@              2@      @                              0@       @              @       @      F@      �?      1@      �?      �?              T@      _@      �?      @     �P@      @      t@      D@      h@     �R@      @              I@     �U@                     �C@      @      j@      4@      `@     �H@      @              A@     �M@                      :@       @     �[@      ,@     @V@     �B@      @              0@      <@                      *@      �?     �X@      @      D@      (@       @              >@     �B@      �?      @      ;@       @     �\@      4@     �O@      9@                      <@     �A@      �?      @      ;@       @     �M@      4@     �@@      7@                       @       @                                     �K@              >@       @              8@      k@     `x@      <@     �I@     �u@     @R@     8�@      g@      @     �p@      :@      @      ,@      P@       @      @      ;@      @     �a@      *@     �P@      5@              @       @      ,@       @      @      (@      @      3@       @      2@      @              @      @      @                      @      @      *@      @      @      @                      @      $@       @      @      @              @      @      (@      �?                      @      I@               @      .@              _@      @     �H@      .@                      @      @@                      &@             @[@      @      C@      *@                              2@               @      @              .@              &@       @              4@     @i@     `t@      :@      G@     �s@     �Q@     �{@     �e@     �z@      o@      :@      .@     �_@     `h@      2@      B@     �l@      K@      f@     �a@     `i@      e@      7@      @     �Z@     �c@      ,@      :@      f@      E@      b@     @X@      f@     @^@      4@      $@      4@     �C@      @      $@      J@      (@      @@     �F@      :@      H@      @      @      S@     ``@       @      $@     @V@      0@     �p@      >@     �l@      T@      @              H@      [@      @      @      D@      (@      j@      ,@     �c@     �K@       @      @      <@      7@       @      @     �H@      @      L@      0@     @Q@      9@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @À�uHd@�	           ��@       	                    �?���0��@�           ��@                           �?���j��@�           h�@                          �8@�h��3@�            ps@������������������������       ����>B�@�             m@������������������������       ��v��:@5            �S@                           �?����@�            `u@������������������������       �T�v,Z@�            �o@������������������������       ���x�� @=            �V@
                           �?
�.s�	@�           �@                           �?M���?�	@�           ��@������������������������       ����@           0}@������������������������       ��,
@�           ��@                            @B����@�            �y@������������������������       �R`�FP@�            �q@������������������������       ��Q6�1@P             `@                           �?���@           �@                            �?�%�0@[           ��@                           �?m�+���?L             \@������������������������       �[��⼩�?&            �L@������������������������       �8�+��� @&            �K@                           �?㭫�v8@           �z@������������������������       �8�Zbo�@�            Pp@������������������������       ����r���?h            @e@                           !@ʊ*���@�           p�@                           �?M�l�@�           0�@������������������������       �~�[�s@*            �Q@������������������������       ��J`1J@�           �@������������������������       ��J�'~x�?             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     s@     �@     �B@      M@      }@     �U@     @�@     �j@     X�@     `u@     �@@      ,@      l@     �t@      <@      G@      u@     �P@      y@      f@     �v@      n@      =@              Q@     @U@      �?      @     �T@      $@     @f@      3@     @b@     �K@      @              6@     �B@      �?      @     �E@      "@     @X@      ,@      K@      >@                      &@      <@      �?      @      <@      @     �V@      "@     �C@      1@                      &@      "@              �?      .@      @      @      @      .@      *@                      G@      H@              �?      D@      �?     @T@      @      W@      9@      @             �B@      G@              �?      B@             �E@      @      O@      5@       @              "@       @                      @      �?      C@      �?      >@      @      �?      ,@     �c@     �n@      ;@     �D@     �o@     �L@     �k@     �c@      k@      g@      :@      ,@     @_@     �d@      :@      <@     �g@     �D@     �`@      ]@      e@     `c@      9@       @      =@     �Q@      @      2@     �R@      @     �S@     �C@     �S@      M@      @      (@      X@      X@      5@      $@     �\@      A@      L@     @S@     �V@     @X@      2@              @@     �S@      �?      *@      P@      0@      V@     �D@     �G@      >@      �?              5@     �G@      �?      "@      L@      *@     �J@      7@     �C@      4@      �?              &@      @@              @       @      @     �A@      2@       @      $@               @      T@      k@      "@      (@      `@      3@     ��@      C@     |@     �Y@      @              6@     �L@      @      @      :@      �?     �p@      $@     @a@      .@       @                      $@      @              @      �?     �O@      �?      9@       @                              @                       @              B@              ,@       @                              @      @              @      �?      ;@      �?      &@                              6@     �G@              @      3@             @i@      "@     @\@      *@       @              .@      =@              @      2@             @_@      @      M@      @                      @      2@                      �?             @S@      @     �K@      @       @       @      M@     �c@      @       @     �Y@      2@     �t@      <@     ps@     �U@       @       @      L@     �c@      @       @      Y@      "@     �t@      <@     Ps@     �U@       @       @      @      @              �?      @       @      $@       @      9@      @                      J@     �b@      @      @     @W@      @     Pt@      4@     �q@     �T@       @               @      �?                       @      "@                       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��xhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��i�g=@�	           ��@       	                    @��n���@K           �@                          �?@��:A��@(           ��@                            �?��j�0�@           ��@������������������������       �;M	@           �z@������������������������       �4�S4�|@�             y@                           @2�U�nu@             =@������������������������       �7�FikN@
             2@������������������������       ���q`�@	             &@
                          �4@'Z.z!	@#           X�@                           �?��;�nJ@8           P~@������������������������       �4L����?�            �j@������������������������       ��n�@ !@�            �p@                            @�1f(�I@�            `x@������������������������       ��L��h@�             u@������������������������       �"� :�^@             J@                           �?B��"�g@o           �@                          �;@�+���@�           0�@                           �?�� �T`@            �@������������������������       ��֨ }�@�             k@������������������������       ��2�'�	@�           8�@                            @,���	`	@k            �d@������������������������       ����@I             \@������������������������       ��̀�¬@"             K@                          �7@�i��N@�           p�@                          �1@��>��@*            �@������������������������       ����� @�            �n@������������������������       �!9����@�           ��@                            @�#��y{@�            �s@������������������������       �֦1h@�            �n@������������������������       �p��@-            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �p@     ��@      =@     �J@     �z@      U@      �@      k@     ��@     �v@      C@      @      \@     �q@      *@      1@     @g@     �F@     0~@     �V@     �t@      c@      .@      @      P@     �b@      &@      "@     �]@      >@     `b@     @S@     �a@     �X@      $@      @      K@     @b@      &@      "@     @\@      =@     `b@     �R@     `a@     �W@      $@       @      =@     @U@      �?      @     �J@      $@     �R@      K@     �N@     �H@      @       @      9@     �N@      $@      @      N@      3@     @R@      4@     �S@      G@      @       @      $@      @                      @      �?              @       @      @               @      @      @                      @                       @      �?       @                      @                               @      �?              �?      �?      �?                      H@     �`@       @       @      Q@      .@      u@      *@      h@      K@      @              6@     �M@      �?      @      6@      �?      m@      @     �\@      8@                      @      5@               @      @             �_@      �?      G@      @                      .@      C@      �?       @      1@      �?     @Z@      @      Q@      2@                      :@     �R@      �?      @      G@      ,@      Z@      @     �S@      >@      @              :@     �Q@      �?       @     �E@      ,@      U@      @     �O@      9@      @                      @               @      @              4@       @      .@      @               @     �c@     0t@      0@      B@     `n@     �C@     �@     �_@     p~@      j@      7@       @     �V@     �`@      (@      7@     �b@      0@     �b@      U@     �g@      ^@      3@      @     �S@     �]@      "@      ,@     �`@      $@     �`@     �N@     �e@     �S@      .@              5@     �A@                      6@             �I@      @      O@      1@      @      @     �L@      U@      "@      ,@      \@      $@      U@     �K@     �[@     �N@      (@      �?      *@      *@      @      "@      1@      @      0@      7@      3@      E@      @      �?      "@      @      �?      @      *@      @      "@      ,@      1@      ?@      @              @      $@       @      @      @      �?      @      "@       @      &@      �?             �P@     �g@      @      *@      W@      7@     `v@     �E@     �r@     @V@      @              D@     @c@      @       @     �K@      &@     �r@      0@     �k@      K@      @              @      @@                       @             �X@      @      U@      $@       @              B@     �^@      @       @     �G@      &@     �i@      $@      a@      F@      �?              ;@     �B@              @     �B@      (@     �K@      ;@      S@     �A@      �?              *@      @@              @      @@      (@      C@      6@     �O@      =@      �?              ,@      @              �?      @              1@      @      *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ꤂ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��זw@�	           ��@       	                   �1@Al��$�@F           Ҡ@                            �?��w[+r@�           P�@                           �?�Q�V-;@c            �c@������������������������       ��mr��@!             L@������������������������       ������?B            @Y@                           @��ے$@           �|@������������������������       ����c�@�            `j@������������������������       ����Hk@�            @o@
                          �4@j�C��@�           ��@                           �?b��v@�            �@������������������������       ��C���@�             x@������������������������       ����\=�@�           @�@                            �?[A�{@@�            pw@������������������������       �睁��@~            �i@������������������������       �n뮗<�@m            @e@                          �;@����@N           ��@                           �?ͥ�Oj@:           ��@                          �:@����T@�            �v@������������������������       �d����`@�            �s@������������������������       ���B@�U @             H@                           @a�˵'	@^           �@������������������������       ��aU��	@y           ؂@������������������������       �w��7?@�            �v@                           @�NYtE	@           P{@                           @rYw�<�	@�             t@������������������������       ��q�|	@}            �i@������������������������       ��j��q�@O            �]@                          �=@��Z�Ai@H            �\@������������������������       ��ґ�h@(            @Q@������������������������       ���	���@              G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     �o@     ȁ@      :@      L@     �}@     �V@     (�@      l@     Ȉ@     0v@     �E@      "@     �X@     �s@      *@      .@     �l@      D@     P�@     �V@     ~@     @d@      2@       @      9@     �U@       @       @     �G@      @     �p@      7@     �]@     �B@      @              @      5@              �?      *@      @     �R@       @      0@      0@                      @      $@                      $@      @      *@      @       @      @                              &@              �?      @             �N@      @       @      *@               @      5@     @P@       @      �?      A@             @h@      .@     �Y@      5@      @              *@      0@                      .@             �[@      $@     �B@      @      @       @       @     �H@       @      �?      3@              U@      @     �P@      ,@              @     @R@     �l@      &@      *@     �f@      B@     �y@      Q@     �v@     @_@      .@      @     �N@     �c@       @      (@     �`@      2@     pt@     �J@     �p@     @Z@      (@              0@      E@               @      7@      �?     �d@      $@     @X@      ;@       @      @     �F@     @]@       @      $@     �[@      1@     `d@     �E@     @e@     �S@      $@       @      (@     �Q@      @      �?     �H@      2@     �U@      .@     �W@      4@      @      �?      @     �I@       @      �?      0@      .@      B@      &@     �N@      @      �?      �?      @      3@      �?             �@@      @     �I@      @      A@      .@       @      2@     �c@     �o@      *@     �D@      o@      I@     �s@     �`@     �s@      h@      9@      @     �_@     @g@      "@      @@      g@      =@     pp@     �Z@     �o@      [@      4@             �A@      L@      �?      @     �@@              Y@      .@     �V@      :@                      A@     �D@      �?      @      >@             @T@      .@     �T@      8@                      �?      .@                      @              3@               @       @              @     �V@     @`@       @      <@      c@      =@     `d@      W@     @d@     �T@      4@      @     �Q@      U@      @      4@     @Y@      3@      Q@     �R@     �U@      K@      1@      �?      5@      G@      @       @     �I@      $@     �W@      2@      S@      <@      @      (@      ?@      Q@      @      "@      P@      5@      J@      :@      N@     @U@      @      (@      7@     �H@      @      @     �H@      4@      <@      9@      @@      Q@      @      &@      (@      =@      �?      @      =@      .@      5@      ,@      .@      H@       @      �?      &@      4@      @              4@      @      @      &@      1@      4@      @               @      3@               @      .@      �?      8@      �?      <@      1@                      @      2@                      @              3@              2@      @                      @      �?               @      "@      �?      @      �?      $@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJP�MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�k�ѨR@�	           ��@       	                    �?�e��^�@l           �@                          �8@�\x�@�           ؃@                           �?E0J�B@4            }@������������������������       ��`6@�             t@������������������������       ���5=52@W            @b@                            �?�SN�@k             e@������������������������       ��Z��<@5            @U@������������������������       �Zz�eF@6             U@
                           �?U|��Fv	@�           �@                           @�N���	@�           x�@������������������������       �u��:�[	@w           ��@������������������������       �Թ��F�	@R             a@                          �1@��+�=�@           �z@������������������������       ��&��>@'            �O@������������������������       ����ܥ@�            �v@                           @%����@7            �@                          �1@Re�-��@'           �@                           @�]�t�?�            �j@������������������������       ���R�c0�?5            �U@������������������������       �G��i���?O            �_@                           @��aaJ@�           X�@������������������������       ��VM@v           ��@������������������������       ��,�8��@-            @S@                           @Sa�I\@           8�@                          �5@�x�	@�            �t@������������������������       ���4�] @�            �k@������������������������       �j����@:            @[@                            �?��/f�@H           �@������������������������       �E��7@�            �r@������������������������       �ʜ�[@�             j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     �p@     ��@      7@     �N@      ~@     �P@     8�@     �l@     8�@     v@      C@      ;@     �h@     �t@      1@     �F@     �t@     �K@     �t@     �g@      x@     �m@      ?@      �?     �L@     �V@       @      &@     @S@      @      c@     �B@     `b@     �I@      @             �E@      P@       @      @     �G@      �?     �`@      5@      ^@      =@      �?             �A@     �I@       @      @     �A@      �?     @R@      4@      T@      3@      �?               @      *@               @      (@              N@      �?      D@      $@              �?      ,@      :@              @      >@      @      4@      0@      ;@      6@      @      �?      @      1@              �?      @       @      @       @      .@      1@      @              @      "@              @      7@       @      *@       @      (@      @              :@     `a@      n@      .@      A@      p@      I@     @f@      c@     �m@      g@      ;@      :@      ]@      f@      .@      6@     �g@      A@     �W@     �Y@     �e@     �a@      9@      4@      Y@     �c@      *@      6@     @e@      ?@     �U@     @S@     �c@     @`@      *@      @      0@      2@       @              5@      @       @      :@      *@      (@      (@              7@      P@              (@     @P@      0@     �T@     �H@     �P@     �E@       @              @       @                      @              8@      .@      @      @                      2@      L@              (@     �N@      0@     �M@      A@      P@     �C@       @      �?     @Q@     �l@      @      0@     �b@      &@     ��@     �D@     Pz@     @]@      @      �?     �B@      Z@      @             �Q@      @     �w@      5@     �k@     �G@      @              @      "@                      @             �a@       @     �I@      @                      @      @                      �?              M@       @      *@      @                              @                       @             �T@              C@       @              �?      A@     �W@      @              Q@      @     �m@      3@     `e@     �D@      @      �?      <@     @T@      �?             �M@      @     @l@      &@     @d@      ?@                      @      ,@       @              "@      �?      (@       @      "@      $@      @              @@     �_@      @      0@     �S@      @      r@      4@     �h@     �Q@      �?               @     �M@              @      :@             �`@      @     @T@      2@                      @      B@              @      "@             �Y@              L@      (@                      @      7@                      1@              >@      @      9@      @                      8@     �P@      @      (@      J@      @     �c@      1@     �]@      J@      �?              (@     �C@              $@      @@      @      V@      "@     �S@      ;@                      (@      <@      @       @      4@             �Q@       @      D@      9@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��J9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�-J�o@�	           ��@       	                    �?O���@r           x�@                            �?R�m���@           0�@                           @f�^���@$           }@������������������������       �[���?z@�            �r@������������������������       ����ڙ@l             e@                           �?��Y��@�            Py@������������������������       �֛�h�@K            @`@������������������������       ��T���@�            0q@
                           �?�����@T           X�@                           �?�k
~�@�            @w@������������������������       ����@^@�            @q@������������������������       �L���<�@<             X@                           @��5�q	@s           �@������������������������       ��̵��*	@           ��@������������������������       ���G�A�@V            �a@                           @b4e�7�@           4�@                          �1@�i���@�           �@                          �0@��G��5�?�             p@������������������������       �v)`V��?5            @T@������������������������       �P�WAߦ�?i             f@                          �5@:{��@6           ��@������������������������       ����H�@?           �~@������������������������       �Y��W��@�            �x@                          �5@��F��@J           ��@                            @�*Э�@�            �q@������������������������       ��ۚ�+@�            �k@������������������������       �J}�5u��?,            �O@                            �?������@�            �n@������������������������       ����KY�@$             K@������������������������       �a���Ti@p             h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     @r@     x�@      E@      I@     0~@     @T@     (�@     �j@     x�@     pv@      C@      0@     �l@     �s@      ?@      E@     0u@      N@     �w@      f@      w@     �n@      ?@      "@     �S@     ``@      1@      &@     �a@      >@     `d@     �P@      _@      V@      "@      �?      =@     @T@      @      @     @S@      4@      V@     �H@      L@      G@      @      �?      7@      F@      �?      @      L@      "@     @Q@      .@     �D@      ?@       @              @     �B@      @       @      5@      &@      3@      A@      .@      .@      @       @      I@      I@      &@      @     @P@      $@     �R@      2@      Q@      E@      @              1@      *@       @      @      8@      @      B@      �?      3@      "@      �?       @     �@@     �B@      "@             �D@      @     �C@      1@     �H@     �@@       @      @     �b@      g@      ,@      ?@     �h@      >@     `k@     @[@     �n@     �c@      6@              F@     �L@              @      A@             @R@      ,@     @Z@     �A@      @             �A@      I@              @      ?@              F@      $@      Q@      >@      @              "@      @                      @              =@      @     �B@      @       @      @     �Z@      `@      ,@      :@     `d@      >@     @b@     �W@     `a@     �^@      1@      @     �X@     @Z@      ,@      9@     @a@      8@     �^@     @R@     @`@     �[@      @      @       @      7@              �?      9@      @      8@      6@      "@      (@      $@      �?      O@     `n@      &@       @      b@      5@     8�@      B@     �y@     �\@      @      �?      C@     �e@       @      �?     �T@      ,@     �|@      9@     @q@      R@       @              �?      C@                      *@             �a@              L@       @                              6@                                      =@              :@      @                      �?      0@                      *@             @\@              >@      @              �?     �B@     �`@       @      �?     @Q@      ,@     �s@      9@     �k@      P@       @              $@      S@      �?      �?      ;@      &@     �h@      &@     �^@      A@      �?      �?      ;@      M@      �?              E@      @     @^@      ,@     @X@      >@      �?              8@     �Q@      "@      @      O@      @     `c@      &@     `a@      E@      @              @      F@      @      @      <@             �Z@      @      Q@      1@      @              @     �E@      �?      @      9@             @Q@      @     �L@      &@      @               @      �?       @      �?      @             �B@              &@      @                      1@      ;@      @       @      A@      @     �H@       @     �Q@      9@                      "@                              @      @      ,@      @      1@       @                       @      ;@      @       @      <@      @     �A@      @      K@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJZ� hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�k�!8K@�	           ��@       	                    �?��)���@           ��@                          �5@�c�3,@�           ؃@                            �?�m�eѧ@�            �x@������������������������       �`/wp@�@�            �k@������������������������       �#�*��?m            �e@                          �<@n�D*B�@�             n@������������������������       �@�a|�@{            `h@������������������������       �yz�m+@            �F@
                          �=@0%�O$_@s            �@                          �8@���ew�@c           P�@������������������������       �6�0@)           �}@������������������������       ���-hR�@:            �T@                          �?@�4�XK@             :@������������������������       ���qa@	             .@������������������������       ��A5���?             &@                           @G�:$T@�           �@                           @|��,^n	@�           H�@                          �9@A����_	@u           $�@������������������������       ����,�@�           (�@������������������������       �mu,ݚ
@�            �l@                          �:@Xj�i��@G           H�@������������������������       �<��:~[@           �z@������������������������       �L��;x@B            �W@                           @����W@�           ��@                          �1@�	���@	           p�@������������������������       ����@�?b             c@������������������������       �s^N��@�           ��@                          �;@��E�@�            �t@������������������������       ����
�*@�            �q@������������������������       �:.�_|�@              H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     `q@     �@     �G@     �G@     |@     �Q@     `�@     �k@     ��@     �u@      ;@              S@     `e@      @      @      X@       @     p{@      =@     �r@     �T@      @              D@     @S@      @      @     �G@      @     �o@      1@     �`@      H@       @              (@     �G@                      4@      @     `h@      &@      T@      7@       @              @      ?@                      0@      @     @X@      @     �G@      0@       @              "@      0@                      @      �?     �X@      @     �@@      @                      <@      >@      @      @      ;@       @      M@      @     �K@      9@                      8@      0@      @      @      8@      �?      L@      @     �H@      *@                      @      ,@               @      @      �?       @      �?      @      (@                      B@     �W@      �?             �H@      �?     @g@      (@     �d@      A@      �?              B@     @W@      �?             �D@      �?     �f@      @     �d@      ?@      �?              @@      R@      �?              ;@             @e@      @     �a@      7@      �?              @      5@                      ,@      �?      (@              6@       @                              �?                       @              @       @       @      @                              �?                      @              @      @      �?      @                                                      @              �?      @      �?                      8@     @i@     p{@     �E@     �D@     v@      O@     ��@      h@     �~@     `p@      8@      8@      `@     �p@      =@      =@      n@      H@     �h@     `d@      l@     `f@      4@      2@     @V@      e@      8@      3@     `f@      B@      `@     �P@     �d@      `@      (@       @      M@     �`@      $@      0@     �b@      9@     @]@      G@      b@      W@      @      $@      ?@      B@      ,@      @      >@      &@      &@      5@      4@      B@      @      @      D@      Y@      @      $@      O@      (@     �Q@      X@     �N@     �I@       @      @      >@     �X@      @      "@      K@       @      M@     �S@      H@      ;@      @      �?      $@       @              �?       @      @      (@      2@      *@      8@       @             @R@     @e@      ,@      (@      \@      ,@     �v@      =@     �p@     �T@      @              G@      `@       @       @     �R@       @     �r@      1@     �g@     �G@      @              @      ,@                      $@             �S@              B@       @                     �D@     �\@       @       @      P@       @     @k@      1@      c@     �C@      @              ;@      E@      (@      $@      C@      @     �Q@      (@     @S@      B@                      5@     �A@      "@      "@      9@      @     �P@      (@     @R@      ;@                      @      @      @      �?      *@      �?      @              @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���M@�	           ��@       	                    @�`Ar4�@           ��@                          �7@y��(-@�           H�@                          �4@K���}�@           �z@������������������������       ����xk@�            �p@������������������������       �1���Ћ@g             d@                            @Sa`��@�            �k@������������������������       �Ѓz�9@b            �b@������������������������       ��<}O��@,            �Q@
                            @� ���)@]           8�@                           @��v���@            @|@������������������������       �E �7 @�            �s@������������������������       ��vfp@Y            �a@                           @��UÔ�?=            �X@������������������������       ����H�b�?             D@������������������������       ��P\"�'�?%            �M@                           �?�b��h(@�           2�@                            @	�m	@q            �h@                            �?n�m��K	@J            �`@������������������������       ��3�B�	@*            �T@������������������������       �������@              I@                           �?gu���N@'             P@������������������������       ��rh�p�@             5@������������������������       �x�s�:�@            �E@                           @$6�7��@(           ��@                          �8@Nf��b	@�           x�@������������������������       �ca��@�           �@������������������������       �戹�G2
@           �y@                           @�q�ܓ[@�           ؐ@������������������������       �|�YB@�           ��@������������������������       ����>C�@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �p@     �@     �C@     �L@     `~@     @R@     ��@     �m@     �@     `v@      @@              T@     `b@      @      &@     �_@       @     0z@      8@     r@     �T@      @             �O@     �T@       @      $@     @X@      @     �b@      .@     �c@     �N@      @             �D@     �I@               @     �K@      @     �]@      @     @[@     �D@      �?              (@     �B@               @     �B@      �?     �Q@      @     �R@      ;@      �?              =@      ,@                      2@       @     �G@       @      A@      ,@                      6@      ?@       @       @      E@       @      @@      "@      I@      4@      @              0@      5@              @      7@       @      6@      @     �B@      3@      @              @      $@       @      @      3@              $@      @      *@      �?                      1@     @P@      @      �?      >@      @     �p@      "@     @`@      6@                      ,@      P@      @      �?      ;@      @     @j@       @     �X@      6@                      (@      D@                      .@       @     �d@      @     �O@      *@                       @      8@      @      �?      (@      �?      G@      @     �A@      "@                      @      �?                      @             �M@      �?      @@                              �?      �?                                      =@              "@                               @                              @              >@      �?      7@                      ,@      g@     �x@      @@      G@     pv@     @P@     p�@     �j@     �@     0q@      ;@       @      1@      :@              @     �B@      @      1@      4@      A@      6@      @      @      "@      ,@              @      5@      @      0@      @      ?@      .@      @      @       @      &@              �?      ,@      @       @      @      (@      *@      @      @      �?      @               @      @      @       @      �?      3@       @              �?       @      (@                      0@      �?      �?      *@      @      @       @      �?               @                      �?                      @              @       @               @      @                      .@      �?      �?      "@      @       @              @      e@      w@      @@     �E@      t@      M@     �@      h@      ~@     �o@      5@      @     �\@      k@      =@      B@     �j@      L@     @k@     �c@      j@     �d@      1@      @     @T@      b@      &@      <@     @e@      @@      g@     �W@     �c@      ]@      @      @     �@@      R@      2@       @      E@      8@      A@      P@     �J@     �H@      (@              K@     �b@      @      @     �[@       @     0v@     �@@     �p@      V@      @              >@     @\@      �?       @     �R@      �?     0r@      5@      i@     �K@       @              8@      C@       @      @      B@      �?      P@      (@     �Q@     �@@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJwmRhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�����f@�	           ��@       	                     @'��4�@!           ؓ@                          �8@\�=�@S           0�@                           @��l��@�           0�@������������������������       �#_��d@�            @s@������������������������       ���_p@!            }@                            �?E��#�@n             d@������������������������       �pX�+�%@V             _@������������������������       �Ͱ��F5@             B@
                          �2@��"�w@�             u@                           @�Ԇ{Dw@D             ^@������������������������       ��!Ǘm�@&            �M@������������������������       �q���(�?            �N@                          �9@lW�e@�             k@������������������������       ��'�D0@d            @b@������������������������       ��b�@&            �Q@                           @���2@@�           ��@                          �5@H��)��@�           �@                           �?��w��U@            ��@������������������������       �A����8@           �{@������������������������       ����@           `�@                           �?u�M5+	@�           ��@������������������������       �>/k��@>             X@������������������������       ��=i
��@Y            �@                            �?���v0	@�            �t@                          �3@8��f1	@y            `i@������������������������       �����,�@"             K@������������������������       �2j��@W            �b@                          �<@=:���@W            @`@������������������������       ��˲Ctx@N            @\@������������������������       ���a{��?	             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     Ё@      >@      J@     �}@     �V@     x�@     @l@     ��@     v@      @@       @     @U@     @g@      @      (@     �\@      (@      |@     �G@     �p@     �U@      @       @     �M@      b@       @      @     �T@      $@     �t@      >@      i@     �M@      @             �H@     �[@       @      @     �P@      @     `s@      1@      e@     �B@      @              =@      >@      �?      @     �C@      �?     �V@      *@     �T@      .@      @              4@     @T@      �?              ;@      @     �k@      @     �U@      6@               @      $@      A@              �?      1@      @      7@      *@      @@      6@      �?       @      "@      :@              �?      $@      @      1@      *@      4@      4@      �?              �?       @                      @              @              (@       @                      :@     �D@       @      @      ?@       @     �\@      1@      Q@      ;@                      @      @              @      @       @     @P@      @      6@      @                      @      @              @      @       @      6@      @      $@      @                      �?      @                      �?             �E@              (@      �?                      3@      A@       @      @      :@              I@      ,@      G@      6@                      2@      =@       @       @       @              =@       @     �@@      1@                      �?      @              �?      2@              5@      @      *@      @              0@     `j@      x@      :@      D@     `v@     �S@     x�@     `f@     @     �p@      ;@      $@     `e@     �u@      9@     �B@     �s@     �P@     �~@     �`@     �|@      m@      2@      @     �O@      k@      &@      (@     �b@      2@     �t@     �O@      q@     @Z@      @      @      @@      R@      @      @     �Q@      @      Q@      A@     �U@     �I@       @              ?@      b@      @      @     @S@      &@     �p@      =@     `g@      K@      �?      @      [@     @`@      ,@      9@     �d@     �H@      d@     �Q@     �g@      `@      .@       @      ,@      $@              @      ;@       @      @      $@      "@      @      @       @     �W@      ^@      ,@      5@      a@     �D@     �c@     �N@     `f@      _@      $@      @      D@      C@      �?      @      G@      (@      P@     �F@     �A@      A@      "@      @      9@      5@      �?      @      8@      &@      @@     �A@      7@      7@      �?              @      @               @      @      �?      0@      �?       @      *@      �?      @      5@      0@      �?      �?      5@      $@      0@      A@      .@      $@               @      .@      1@                      6@      �?      @@      $@      (@      &@       @      �?      &@      0@                      ,@      �?      @@      $@      "@      &@       @      �?      @      �?                       @                              @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�IchG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��ň'@�	           ��@       	                    �?��MCz@f           �@                           �?�j��@           \�@                           �?l>]�@;           �~@������������������������       �-�#LQ�@z            @h@������������������������       ��4A4A@�            `r@                           @�G��e	@�           ��@������������������������       ��B�B�	@r           ��@������������������������       �����	@T            @_@
                           �?! u1�@e           ��@                          �=@�ȏe�@�             j@������������������������       ���	�%@�            �h@������������������������       ��7���� @             &@                           �?�U�1 �@�            0v@������������������������       �Q��h�@<             U@������������������������       �puy��@�            �p@                           �?�Qg�&@8           ��@                           @	�q�� @\           ��@                           @i��1�?�            �u@������������������������       �	C�o�b @\            �`@������������������������       �����H�?�             k@                           �?Jd�Z�@z            �g@������������������������       ����V�?<            �V@������������������������       �jN9܅�@>            �X@                           @����pC@�           ��@                           @�]�~U@           p�@������������������������       ��ϋ0��@;            �@������������������������       �xz3� @�            �t@                            �?)n�S�O@�            Pu@������������������������       ��5w���@0            @T@������������������������       �-,z?�Z@�            @p@�t�b�     h�h5h8K ��h:��R�(KKKK��h��B�        0@     pr@     ��@      <@     �E@     �~@      S@     h�@     �i@     ��@     �v@     �@@      0@     �h@     t@      .@      ?@     @v@      N@     �u@     �d@      y@     �o@      8@      0@      d@     �l@      .@      <@     �q@      H@     �j@     �_@     �q@     @i@      4@             �E@     @R@      �?       @     @R@      �?     @Y@     �@@      Z@      I@      �?              1@      9@                      >@             �G@       @      K@      (@      �?              :@      H@      �?       @     �E@      �?      K@      9@      I@      C@              0@     @]@     �c@      ,@      4@     �i@     �G@     �\@     @W@     @f@      c@      3@      $@     �Z@     �a@      *@      2@      f@     �C@     @Z@     �T@     `e@     `a@      $@      @      &@      2@      �?       @      ?@       @      "@      $@      @      *@      "@             �B@     �V@              @      S@      (@     �`@     �C@     �]@     �I@      @              *@      ?@              �?      =@      @      H@      .@     �E@      7@      �?              &@      ?@              �?      :@      @      H@      &@     �E@      6@      �?               @                              @      �?              @              �?                      8@     �M@               @     �G@       @     @U@      8@     �R@      <@      @              @      "@                      @      �?      6@      @      ?@      �?      @              1@      I@               @      D@      @     �O@      5@      F@      ;@                     �X@      n@      *@      (@     @a@      0@     ��@     �C@     �x@      [@      "@              6@     �R@      �?       @      ;@      @     �p@      @     �\@      1@       @              0@      E@                       @      @     �h@       @     @Q@      (@                      @      9@                      @             �P@              7@      "@                      "@      1@                      @      @     �`@       @      G@      @                      @     �@@      �?       @      3@              R@      @     �F@      @       @               @      2@               @      @              F@              2@                              @      .@      �?              (@              <@      @      ;@      @       @              S@     �d@      (@      $@     �[@      *@      x@     �@@     �q@     �V@      @             �I@      ]@      @      @     �S@      @     �r@      ,@     �j@      L@      @             �D@      Q@      @       @     �K@      @     �d@      *@     �\@     �E@      @              $@      H@              �?      7@             �`@      �?     @Y@      *@                      9@      I@       @      @     �@@       @     @V@      3@     �P@     �A@                       @      @                      @       @      ?@      &@      (@      @                      1@     �F@       @      @      ;@      @      M@       @     �K@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�5�[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @
u8��e@�	           ��@       	                     �?ƌ�8�@l           4�@                           �?A��f�@�           H�@                           �?�c� @�            x@������������������������       ���5���@�            0q@������������������������       ��J	H�M@E            �[@                           @=�*��	@�           ��@������������������������       �Y���m;	@3           �~@������������������������       ��7�h	@�            pr@
                           �?�FX�,�@�            �@                           �?�B3�@	@�           ��@������������������������       �F-[o��@�             n@������������������������       ��l}uf	@H           �@                            @�~�]G@�            `q@������������������������       �K�fĖ@:            �X@������������������������       �)>����@p            �f@                          �2@�RV�� @#           ��@                           @R�0&z� @Z           �@                          �1@s�+0ʿ�?�            �s@������������������������       ��iҴ�?v            @h@������������������������       ��67^��@I            �]@                          �0@QH���@�            �l@������������������������       �f��	�?              L@������������������������       �u=�I�@{            �e@                           �?�����&@�           H�@                          �>@m�@�             v@������������������������       ����@�             u@������������������������       �      @
             0@                           @´����@�           ��@������������������������       ���.�U�@�           ؈@������������������������       �v�E���@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     pr@     ��@      ;@     @P@     }@     �Y@     ؍@     �k@      �@     `u@      6@      ,@      j@     @u@      4@     �K@     �s@     �U@     `v@     �e@     �w@      m@      3@      @     �Z@     @f@      "@      8@     `a@      M@     `k@     �X@      i@     �]@      ,@      �?     �@@     �I@               @      ;@      �?     �\@      6@     @V@     �@@      @      �?      <@     �E@              @      9@             �O@      4@     �L@      ?@      @              @       @              @       @      �?      J@       @      @@       @       @      @     @R@     �_@      "@      0@      \@     �L@      Z@      S@     �[@     @U@      "@       @     �E@     �U@      @      "@     �Q@      D@      O@      <@      R@      P@      @      @      >@      D@      @      @      E@      1@      E@      H@     �C@      5@       @      @     �Y@     @d@      &@      ?@     �e@      =@     `a@     @S@     �f@     �\@      @      @     �S@     �^@      $@      <@     �`@      5@     �T@      L@     @_@     @U@      @              *@      C@      @      (@     �H@      @     �A@      .@     �G@      8@              @     �P@     @U@      @      0@     �T@      1@      H@     �D@     �S@     �N@      @              8@     �C@      �?      @     �D@       @      L@      5@      L@      =@                      @      @                      7@      @      *@      (@      9@      "@                      2@      A@      �?      @      2@      @     �E@      "@      ?@      4@               @     �U@      l@      @      $@      c@      0@     ��@      H@     p|@     �[@      @              <@     �O@      @       @      5@             �o@      @     �a@      6@                      4@      =@      @               @             �c@      @      U@      @                      "@      "@                      @             @]@              I@      @                      &@      4@      @              @              D@      @      A@      @                       @      A@               @      *@             �X@      �?      M@      .@                              (@                                      8@              (@       @                       @      6@               @      *@             �R@      �?      G@      @               @      M@      d@      @       @     �`@      0@     `u@      F@     �s@      V@      @              @     �M@       @      �?      :@      @     ``@      @     @Z@      *@                      @      M@       @      �?      6@      @     @`@      @     @Y@      "@                              �?                      @      �?      �?      �?      @      @               @     �J@     �Y@      �?      @     �Z@      $@     `j@      D@      j@     �R@      @       @     �I@     @Y@      �?      @     �X@      @     `j@     �A@     �i@      R@      @               @      �?                      @      @              @       @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�LfhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?K1>��x@�	           ��@       	                    �?O���@           T�@                           �?A2��1@8            @                            �?����g@x            �h@������������������������       ��1C�Bf@K            ``@������������������������       ��v	^&�@-            �P@                          �7@�=����@�            �r@������������������������       �����@�            �h@������������������������       ���e@�@>            �X@
                          �4@9��d2P@�           (�@                           @a�ҫi@ @
           `y@������������������������       �
��X@k            �c@������������������������       ���t����?�             o@                          �=@���@�
@�            �t@������������������������       �T�9��G@�            Ps@������������������������       �l�:.1�@             :@                          �5@\�s��l@�           �@                           @�-0���@s           �@                           �?��t�c@�           0�@������������������������       �qW�5��@4           �~@������������������������       �F�'��/@�            �k@                          �4@b�Q��@�           �@������������������������       ����޶@j           H�@������������������������       �eT���@F             ]@                          �<@{�c��	@           ē@                           �?:5�9�K	@~           P�@������������������������       ���6e@�             y@������������������������       �x-�[�	@�           Ђ@                            �?}����z	@�            pp@������������������������       �����sU@O            �a@������������������������       �{�Z���@M            �^@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      s@     P�@      B@     �N@     0~@     �P@     ��@     �m@     ��@     �u@      @@      �?     @W@     �f@      @      @     �^@      $@     �z@      C@     �q@     �Q@       @      �?      J@     �S@       @      @     �T@       @     �V@      9@     �]@     �D@              �?      4@      <@                      ;@             �F@      @      N@      (@              �?      0@      2@                      0@              ;@      �?      D@      (@                      @      $@                      &@              2@      @      4@                              @@      I@       @      @     �K@       @      G@      4@     �M@      =@                      7@     �A@                      =@      �?      C@      $@     �F@      2@                      "@      .@       @      @      :@      �?       @      $@      ,@      &@                     �D@     �Y@       @       @     �D@       @     �t@      *@     �d@      >@       @              9@      G@               @      ,@             @j@      @     �V@      *@                      *@      3@              �?      @              O@       @     �F@      &@                      (@      ;@              �?      "@             �b@      @     �F@       @                      0@     �L@       @              ;@       @     �^@      @      S@      1@       @              ,@      L@       @              7@      @     �\@      @     @R@      0@                       @      �?                      @       @       @      @      @      �?       @      1@     �j@     Py@      @@      L@     �v@      L@     ��@     �h@     0@     0q@      >@      @      P@     �k@      (@      5@     �f@      1@     `w@     �T@     0s@     �\@      &@      @     �C@     �[@       @      1@      ^@      (@     �_@     �P@      _@     @R@      @      @      =@      R@      @      (@     �V@      $@      P@      E@      V@     �N@      @              $@     �C@      �?      @      =@       @      O@      9@      B@      (@                      9@     �[@      @      @      N@      @      o@      0@     �f@     �D@      @              8@     @W@      @      @      H@      @      j@      0@     �b@      C@                      �?      1@              �?      (@       @      D@             �A@      @      @      $@     �b@      g@      4@     �A@     �f@     �C@      d@      ]@      h@      d@      3@      "@     @\@     �c@      .@      3@     �`@      =@     �a@      U@      d@     �]@      1@      �?      F@     �O@       @      @     �K@      @     �N@      =@      O@      O@      "@       @     @Q@      X@      @      0@      T@      :@     �T@     �K@     �X@      L@       @      �?      B@      9@      @      0@     �F@      $@      1@      @@      ?@     �E@       @              1@      (@              @      1@      @      "@      =@      2@      :@       @      �?      3@      *@      @      $@      <@      @       @      @      *@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�F�QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @i�8S�o@�	           ��@       	                   �4@a�y��@u           z�@                           �?.��(�@'           ��@                           �?�5D߬@�            0s@������������������������       ��BU���@4            @W@������������������������       �3����@�            �j@                          �3@��		�@p           �@������������������������       ��kC�9@           P{@������������������������       �*o�o�@Z             a@
                           �?ˣؚ�	@N           4�@                            �?�'BLT�@�            �x@������������������������       ���L��R@�            �k@������������������������       �p�+���@l             f@                           �?P�"��	@[            �@������������������������       ����st>
@�           �@������������������������       �oG����@�            �k@                           �?њ7y7@           0�@                           �?�)��	@a           H�@                            �?4�ʻ@�            `t@������������������������       ���^;�<�?$             O@������������������������       �,�:;\@�            �p@                          �2@�N��� @�            0p@������������������������       ��V�ޟ��?>             Z@������������������������       ��zE�۠ @X            `c@                           @�i@�H\@�           �@                          �7@�:�r�3@�           �@������������������������       ���z��@           ��@������������������������       ���m� @l            `e@                           @���$@�             t@������������������������       �)�.�b5	@+             P@������������������������       ��E�Tr�@�             p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �p@     �@     �A@     �M@     �z@     �T@     (�@      m@     ��@     Px@      <@      4@     �g@     �u@      =@      E@      r@      M@     �w@     `i@     x@      q@      6@      @     �H@     �^@      @      @      Z@      "@      k@     @Q@      i@     @V@      @              .@      G@                      :@      �?     �X@      @     �U@      9@       @              @      3@                      @              >@              ;@      &@                      (@      ;@                      7@      �?      Q@      @      N@      ,@       @      @      A@     @S@      @      @     �S@       @     �]@      O@     @\@      P@      @      @      7@     �O@      �?      @     �I@      @      Z@     �H@     @T@     �H@      @       @      &@      ,@      @              ;@      �?      ,@      *@      @@      .@      �?      .@     �a@      l@      6@     �C@     @g@     �H@      d@     �`@      g@      g@      0@              G@      J@      @      $@      K@      @     @R@      8@      S@      I@      @              6@      8@       @      @      7@      @     �B@      (@     �G@     �B@      @              8@      <@      �?      @      ?@              B@      (@      =@      *@              .@      X@     �e@      3@      =@     �`@      F@     �U@     �[@     @[@     �`@      (@      .@     �R@     �_@      3@      7@     @Z@      C@      O@     �T@      R@     @[@      (@              5@     �F@              @      ;@      @      9@      <@     �B@      :@              @     �R@      m@      @      1@     �`@      9@     h�@      >@     �{@     �\@      @              4@     �V@              �?      9@      "@     Pq@      @     @a@      2@      @              .@     �I@              �?      .@      @      d@      �?      P@      (@                              @                      @      @      C@              &@      @                      .@      H@              �?      (@      @     �^@      �?     �J@       @                      @     �C@                      $@       @     @]@      @     �R@      @      @              @      @                      @             �P@       @      2@              @               @      @@                      @       @     �I@      �?      L@      @              @     �K@     �a@      @      0@     �[@      0@     �s@      :@     s@     @X@      @      @     �C@      [@      �?      @     �R@      @     @o@      *@     �j@     �K@       @              8@     @W@      �?      �?      E@      @     @j@      @     �e@     �D@       @      @      .@      .@              @      @@              D@      @     �D@      ,@                      0@      A@      @      &@      B@      "@      O@      *@     �V@      E@      �?               @       @      @       @      @      @      &@      "@      $@      @                      ,@      :@      �?      "@      >@      @     �I@      @     @T@      B@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ^��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����T@�	           ��@       	                   �<@BR��]F@           h�@                          �1@x���p�@�           �@                          �0@h12��?�            `m@������������������������       ��~�$��?7            �T@������������������������       �
����p�?f             c@                           �?��*p@B           Ȍ@������������������������       �8ĵV�@�            �v@������������������������       �.��؏�@]           p�@
                           �?�퍯6o@6            �U@                           @
,h�{;@            �H@������������������������       �q��5�@             B@������������������������       �g��o��?             *@                          �@@��;�@            �B@������������������������       �J�lf�#@             <@������������������������       �����Z@             "@                          �4@�W�G�Q@�           ޤ@                            �?�QI@�           P�@                           @��?,m�@�            @r@������������������������       ��O��T�@y             g@������������������������       �ޯݩ�{@F            �Z@                          �1@�s�O @           ��@������������������������       �k�8��@�            �o@������������������������       �o����@r           ��@                          �7@��NgV	@�           l�@                           @w֕�.b@�           ��@������������������������       �^��Q��@�            @t@������������������������       ���;P�@�            u@                           �?y�9��	@'           0�@������������������������       ���7�W
@           �|@������������������������       ��Ax��@	           �{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        "@     @s@      �@      ?@     �L@     �{@     �U@     �@     `k@     �@      x@     �A@             �S@     �d@      @      "@     @Y@      @     �}@      H@     @p@     �X@       @             �R@     �c@      @      @     �W@      @     �|@     �C@     �o@     �P@      �?              &@      @@                      ,@              _@       @     �F@      @                       @      .@                      @             �C@              2@      @                      "@      1@                      "@             @U@       @      ;@      @                     �O@      _@      @      @      T@      @     �t@     �B@     �i@     �M@      �?              @@      N@      @      @      C@       @     @R@      =@     @U@      B@      �?              ?@      P@              @      E@      @     Pp@       @     �^@      7@                      @       @              @      @              ,@      "@       @      @@      �?               @      @               @      @              (@      @      @      2@                       @      @               @      @               @      @      �?      2@                                                                      $@              @                               @      @              �?      @               @      @      @      ,@      �?              �?      @                      �?               @      @      @      *@      �?              �?       @              �?      @                      �?              �?              "@     �l@     �w@      ;@      H@     �u@      T@     P�@     `e@     �@     �q@     �@@      �?     �O@     �c@      @      *@     �]@      (@     �t@     �K@     �m@     �Z@      @              1@      @@              �?     �D@      @     @Y@      2@      H@      :@      @               @      0@                      ?@              N@      *@     �@@      7@      �?              "@      0@              �?      $@      @     �D@      @      .@      @       @      �?      G@     �_@      @      (@     @S@      @     �l@     �B@     �g@      T@      @      �?       @      D@      �?      �?      &@              X@       @     �P@      6@                      C@     �U@      @      &@     �P@      @     �`@      =@      _@      M@      @       @     �d@     �k@      6@     �A@     @l@      Q@     �k@      ]@     �p@     �f@      :@       @     �P@      [@      @      6@      X@      .@     @]@      :@     @`@      N@      &@              >@      H@      @      $@     �G@      @      P@      0@     �P@      ?@               @     �B@      N@      �?      (@     �H@      "@     �J@      $@      P@      =@      &@      @      Y@     �\@      .@      *@     @`@     �J@     @Z@     �V@     �a@      ^@      .@      @     �O@     �L@      (@      @      M@      C@     �A@     �N@     �F@      O@      ,@      �?     �B@     �L@      @      @      R@      .@     �Q@      =@      X@      M@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�.�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?<5��}@�	           ��@       	                     @�g?�@           P�@                            �?,$�d��@H           (�@                           �?�$ΞO@�           ��@������������������������       ��K�hl@�            �u@������������������������       ��'*D�X@�            @u@                           @s��4�+@�            �n@������������������������       ��z��z@}            �h@������������������������       ��exBr@             H@
                           �?�Q#.v�@�            �r@                          �1@h�o���@`            �b@������������������������       �TTH&5��?             @@������������������������       �~��Z��@P            @]@                          �3@i[�N�@`            @c@������������������������       �������@.            @S@������������������������       ��Q'~n@2            @S@                          �5@;э�T@�           �@                           �?�:�F�@x           Е@                          �3@ ��5	@A           �@������������������������       ����V�@�            �r@������������������������       �b�X�@�            �j@                           @�Qb��@7           ��@������������������������       ��a�-"T@�            0x@������������������������       ����?��@;           0@                           @��W�R	@!           �@                          �8@��z�	@           ��@������������������������       �kd3ƻ	@�            �v@������������������������       ���`'��	@*           `~@                          �7@��h=^@           �z@������������������������       ����k�@^            @d@������������������������       ��A��@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      s@     �@      ;@     �K@     P}@      X@     �@     �l@     ��@     `w@      >@      �?     �U@     �d@      �?      &@     @]@      3@     p{@     �H@     �p@     �S@      @      �?      M@     �^@      �?      "@      U@      1@     0u@      >@     �i@     �O@      @      �?     �E@     �V@      �?      "@     �P@      (@     �m@      8@     �b@      J@      @      �?      4@      A@      �?       @     �C@      "@     �a@      0@      I@      9@       @              7@     �L@              �?      ;@      @     �W@       @     �X@      ;@      �?              .@      @@                      2@      @     �Y@      @     �K@      &@      �?              ,@      .@                      2@      @     �V@      @      G@      @                      �?      1@                                      (@      @      "@      @      �?              =@     �D@               @     �@@       @      Y@      3@      O@      .@                      &@      .@               @      2@       @     �K@      "@      >@      @                      �?      @                                      2@      @      �?      �?                      $@      $@               @      2@       @     �B@      @      =@      @                      2@      :@                      .@             �F@      $@      @@       @                       @       @                      @              6@       @      ;@      @                      $@      2@                      $@              7@       @      @      @              2@     `k@     �w@      :@      F@      v@     @S@     X�@     �f@     P@     �r@      :@      @     @U@     @i@      "@      3@     @d@      @@     �v@     �Q@     �r@     @a@      "@      @      H@      N@      @      $@     �V@      2@      U@     �D@     �S@     �M@       @      �?      ?@     �@@      @       @      E@      (@     �M@      >@      F@      A@      @      @      1@      ;@       @       @     �H@      @      9@      &@     �A@      9@      @             �B@     �a@       @      "@     �Q@      ,@     Pq@      >@      l@     �S@      �?              4@     @S@              @     �@@      ,@     �Y@      4@     @S@     �B@      �?              1@     @P@       @      @      C@             �e@      $@     `b@      E@              *@     �`@     �f@      1@      9@     �g@     �F@     @h@     �[@     �h@     �c@      1@      (@     @Y@     �_@      0@      2@     ``@      E@      V@     �V@     �W@     �\@      .@      @     �J@      I@      @      .@     �Q@      3@      A@      :@      H@     �A@      @      "@      H@     @S@      $@      @     �N@      7@      K@     @P@     �G@      T@      "@      �?     �@@     �J@      �?      @     �M@      @     �Z@      3@     �Y@     �E@       @              .@      ?@      �?              2@      �?      I@      @      @@      $@              �?      2@      6@              @     �D@       @      L@      .@     �Q@     �@@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��0mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��]�l@@�	           ��@       	                    �?%o-|yK@�           Ԓ@                           �?⹤��@/            ~@                          �1@M����@�            �k@������������������������       �Ή���	�?             ?@������������������������       �g[X���@~            �g@                            @'�"�3@�             p@������������������������       �a��@b             d@������������������������       �zF���@<            �X@
                            �?H�`���@�           ��@                          �9@D�aqM�@r            @g@������������������������       ����"���?f            `d@������������������������       �ۙ>MK@             7@                           @��/*��@\           ؀@������������������������       �?��@A            @Y@������������������������       �T8\I~0@           `{@                          �8@�. �-@�           (�@                           @�a~�B@�           h�@                          �3@~k&��@�           H�@������������������������       ��C��@            �|@������������������������       ��&��@�           P�@                           @��	��~@@           @�@������������������������       ��r�Z9@5           ��@������������������������       �+Kw��)@             1@                          @A@n$M�Ĵ	@�           Ѕ@                          �<@޲��vn	@�           P�@������������������������       ������6	@1           �|@������������������������       ��7���@�             l@������������������������       �|R��>@
             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �q@     �@      C@      N@     �@      V@     <�@      k@     p�@     �u@      2@             @S@     �b@      �?      @      _@      $@      |@     �C@     pp@     �T@      @              G@     �O@      �?      @     �Q@       @      \@      =@     @Y@     �H@      @              5@      =@      �?      @      @@       @     �G@      5@     �C@      9@       @                      @                      @              4@      �?      �?       @                      5@      9@      �?      @      =@       @      ;@      4@      C@      7@       @              9@      A@              �?      C@             @P@       @      O@      8@      �?              .@      .@              �?      =@             �A@      @     �F@      .@      �?              $@      3@                      "@              >@      @      1@      "@                      ?@     �U@              �?      K@       @      u@      $@     @d@      A@      @              �?      5@                      ,@      @     �U@      @      G@      @       @              �?      5@                      (@       @      S@              F@      @                                                       @      @      $@      @       @               @              >@     @P@              �?      D@       @     @o@      @      ]@      ;@      �?              &@      @                      1@      �?      G@      @      *@      @                      3@      O@              �?      7@      �?     �i@      @     �Y@      4@      �?      2@     �i@     �v@     �B@     �K@     Px@     �S@     x�@     @f@     8�@     `p@      (@      (@     `b@     �q@      .@     �B@     @q@     �J@     �@      Z@     �y@      d@      @      &@      V@     �e@      "@      >@      g@     �@@      g@     �V@     �h@     @Y@      @      @      >@     �O@       @       @     @P@      "@     �\@     �A@     @R@      I@       @      @      M@     @[@      @      6@      ^@      8@     �Q@      L@      _@     �I@       @      �?     �M@      [@      @      @     �V@      4@     Pt@      *@     �j@      N@              �?     �L@     �Z@      @      @      V@      1@     Pt@      *@     `j@      M@                       @      �?      �?       @      @      @                      @       @              @      M@      U@      6@      2@     @\@      9@     @T@     �R@      [@     @Y@       @      @     �L@     �T@      2@      2@      \@      6@     @T@     �R@      [@     �X@       @      @     �A@     �L@      *@       @     �O@      &@     �L@      K@     �V@     �M@      @              6@      9@      @      $@     �H@      &@      8@      4@      2@      D@      �?      @      �?       @      @              �?      @                               @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�x�ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?5����@@�	           ��@       	                     �?�9<��@!           ��@                          �;@�^��%@�            �u@                           @�"G�Xv@�            �s@������������������������       �z�f���@{             j@������������������������       ����J���?G             [@                          �=@�l��J	@             A@������������������������       ��}ZG�@             6@������������������������       �^�z|�X@             (@
                           @�m@�o�@K           H�@                          �<@�t����@,           `}@������������������������       �փ��)@           �y@������������������������       �2H�ԗ�@'             L@                           @�G��� @           0{@������������������������       �NH�G#��?�            0r@������������������������       ��,鄘D@_             b@                           @�Y���Y@�           ¤@                           �?o=��	@�           d�@                            �?�N&:n�	@�           ��@������������������������       �j�3�n	@�            �t@������������������������       ��w��	@�            �@                          �5@���J�@�            �v@������������������������       �Ul�>�@�            @j@������������������������       ��h޶�x@g            @c@                          �5@v'��T@�            �@                          �4@����Zc@�           ��@������������������������       �c;,E�@a           �@������������������������       ��B��]q@I             _@                          �<@�L�
��@.           �~@������������������������       ���ղ�@           Py@������������������������       �9Y��P@,             U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     ps@     @�@      @@     �L@     �{@     �P@     �@     @k@     ��@     �v@      9@      @     �U@     `c@      �?      @     �Z@      @     `}@      A@     s@     �S@      @      @      1@     �G@              @      <@       @     �a@      @     �U@      0@      �?              *@      F@              @      :@              a@      �?     �T@      &@                      *@      A@              @      4@             @R@      �?     �L@      @                              $@                      @             �O@              9@      @              @      @      @                       @       @      @       @      @      @      �?      @      @      @                      �?       @      @              @      �?                                                      �?               @       @       @      @      �?             �Q@      [@      �?      �?     �S@      @     �t@      ?@     @k@     �O@       @              J@     �H@      �?      �?     �M@      @     �_@      :@      Z@      H@      �?              G@      E@      �?              H@      @     �^@      .@     @X@     �C@      �?              @      @              �?      &@              @      &@      @      "@                      2@     �M@                      3@       @     @i@      @     �\@      .@      �?              .@      >@                      "@       @     �c@      �?     �P@      "@                      @      =@                      $@              F@      @     �G@      @      �?      8@      l@     �v@      ?@      J@     @u@     �M@     p�@      g@      �@     �q@      6@      8@     �b@     `j@      5@     �C@     `l@      F@     @j@     �c@     @j@     `g@      2@      8@     �^@     �b@      4@      =@     �f@     �A@      a@      `@     @b@      b@      1@      �?      :@      =@      @      $@     �K@      $@     �F@      K@      G@     �C@       @      7@      X@     �^@      ,@      3@     �_@      9@     �V@     �R@      Y@     @Z@      "@              ;@      N@      �?      $@      G@      "@     �R@      =@      P@     �E@      �?               @      C@      �?      @      <@       @      L@      3@      B@      8@                      9@      6@              @      2@      @      2@      $@      <@      3@      �?             �R@     @c@      $@      *@     @\@      .@     �u@      ;@     �r@     �X@      @              6@     @W@      @       @     �E@      @     �n@      $@     `g@      I@      @              6@     �S@      @       @      =@      �?     �j@      "@     @a@      F@                              ,@                      ,@      @     �@@      �?     �H@      @      @             �J@     �N@      @      @     �Q@      $@     @Y@      1@     �\@     �H@      �?             �A@     �I@      @      @      I@      $@     �W@      1@     �Y@      B@      �?              2@      $@      @              4@              @              *@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ
�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�G��9s@�	           ��@       	                   �<@�n�i�@�           t�@                            @�B�_�@�           �@                          �7@Q0�aq�@           ��@������������������������       �4�>PA�@�           �@������������������������       �7��_�@d            `f@                           @��q{��@�            pq@������������������������       �f��Nq@~            �h@������������������������       ���Mv��?0            �T@
                           �?P��@3            �U@                            �?�rsJz@             >@������������������������       �騼����?	             ,@������������������������       �����@
             0@                          �>@4x_�W`@              L@������������������������       �j�w��@             :@������������������������       ��in=��@             >@                           @I\yn�m@�           ؤ@                           @����V@�           r�@                          �1@#���yH	@Y           `�@������������������������       ��z��'@g            �d@������������������������       ���#��	@�           Ȓ@                          �1@�Ѱ&@{           �@������������������������       ���e� @�            @i@������������������������       ���R�@�           ��@                           @����+
@�            0s@                          �:@E�;���	@o            �e@������������������������       �%��1��@T            @_@������������������������       �cnN��;@            �H@                           @�T��@S            �`@������������������������       ���Ƨ@?            @Y@������������������������       �1�0�@             @@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �q@     �@     �@@      M@     �}@     �U@     @�@      l@     ��@     �u@     �D@       @     @U@     `b@      @      $@     @[@      @     �|@     �D@      r@     �T@       @       @     �R@      a@      @      "@     �X@      @     @|@      >@     �q@     �M@      @       @     �I@     �[@       @       @      R@      @     �u@      9@     `j@     �F@      @              C@     �S@       @      �?     �M@      �?     �r@      2@     �d@      ?@      @       @      *@      @@              �?      *@      @     �E@      @     �F@      ,@      @              7@      :@       @      @      :@      �?     �Z@      @     @Q@      ,@                      5@      :@       @      @      5@      �?      K@      @      J@      &@                       @                      @      @              J@              1@      @                      &@      $@              �?      &@               @      &@      $@      7@      �?              �?      @              �?      �?              @      @      @      &@                               @                                      �?      @               @                      �?      @              �?      �?              @              @      @                      $@      @                      $@              @       @      @      (@      �?              @       @                      �?              @       @      @      @      �?              @      @                      "@                      @       @      @              7@     �h@     `v@      =@      H@     �v@     �S@      �@     �f@     �@     �p@     �@@      *@     �d@     �s@      9@      F@     �s@     �Q@     ��@     �b@     �}@     `m@      3@      *@      \@      i@      2@      >@      k@     �J@     `j@     �^@      k@     �c@      2@              @      =@      �?       @      $@              O@      2@      =@      $@              *@     �Z@     �e@      1@      <@     �i@     �J@     �b@     @Z@     `g@     @b@      2@             �K@     @]@      @      ,@      Y@      1@     t@      9@     p@     �S@      �?              @      4@               @      (@             �W@      @     �L@      @                     �H@     @X@      @      (@      V@      1@     `l@      5@      i@      R@      �?      $@      ?@      D@      @      @      G@      "@      H@     �A@     �@@     �@@      ,@      $@      4@      9@      �?       @      B@       @      (@      ;@      "@      .@      "@      @      3@      5@      �?       @      ?@      @      "@      *@      @      "@      @      @      �?      @                      @      @      @      ,@      @      @       @              &@      .@      @       @      $@      �?      B@       @      8@      2@      @              @      (@      �?               @              B@       @      2@      0@       @              @      @       @       @       @      �?              @      @       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJy*3ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�֫��}@�	           ��@       	                    �?
9\�@`           ��@                           �?���,n@�           ��@                           �?���S�@�            �o@������������������������       ��3�&�@I            �]@������������������������       �C���F@S            �`@                          �3@����+� @B           �@������������������������       �9P�����?�            pu@������������������������       �,�P_�*@`            �d@
                            @%#�K,�@�           ��@                           @��w�k	@�           Џ@������������������������       �\^S�K�@"           |@������������������������       ��Y��m@r           ȁ@                           @��2�*w@�            Px@������������������������       �r9��p!@�            �v@������������������������       ��X��\<@             <@                          �<@~�S��@Z           8�@                           �?�î�u@�           \�@                           �?���V�	@�            �@������������������������       �;�i��l	@�            pp@������������������������       �3��J	@           �y@                           @�6��]@�           ��@������������������������       �B��%�@�           Є@������������������������       ��ϲ��[@2            @W@                           @���>�	@�            ps@                          �=@MxT
@�            �m@������������������������       �yAleq&@+            �P@������������������������       �w����$
@o            @e@                           @�c�4��@0            �R@������������������������       �^3
O@             <@������������������������       ��Y�@             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �s@     @�@      <@     �J@     0{@     @U@     ��@      n@     0�@     �v@      B@      @     �\@     `s@       @      ?@     `j@      >@     ��@      W@      @      e@      *@              B@     �Y@       @       @     �J@      $@      t@      4@     @e@      D@       @              0@      C@       @      @      7@      @     �P@      0@     �L@      :@                      @      *@       @              ,@      @     �B@      (@      4@      @                      "@      9@              @      "@              =@      @     �B@      3@                      4@     @P@              @      >@      @     �o@      @     @\@      ,@       @              ,@     �A@              �?      ,@              f@      @      V@      $@       @              @      >@              @      0@      @     �S@      �?      9@      @              @     �S@     �i@      @      7@     �c@      4@     w@      R@     �t@      `@      &@              J@     �a@      �?      2@      Z@      1@     �r@      J@     �l@     �W@      @             �A@     �P@      �?      $@     @Q@      (@     @W@     �D@     �Q@      G@      @              1@     �R@               @     �A@      @      j@      &@     �c@     �H@      @      @      ;@     @P@      @      @      K@      @     �P@      4@      Y@     �@@      @      @      ;@      O@      @      @     �G@      @     �P@      1@     �W@      <@       @       @              @                      @                      @      @      @       @      0@      i@     @n@      4@      6@      l@     �K@     @r@     �b@     @s@      h@      7@      (@     �d@     @j@      *@      0@     �e@     �B@     �p@     �[@     q@     @a@      1@      &@     �W@      ^@      @      &@     @X@      5@     �P@     �Q@      U@     @R@      0@       @     �@@      I@       @      @     �B@      (@      9@      7@      =@      B@      &@      "@      O@     �Q@      @       @      N@      "@     �D@      H@     �K@     �B@      @      �?     �Q@     �V@      @      @      S@      0@     �h@      D@     �g@     @P@      �?      �?      K@     �S@       @      @     �P@      (@     `f@      ;@      f@     �O@      �?              1@      (@      @              "@      @      4@      *@      (@       @              @      A@      @@      @      @     �I@      2@      ;@     �B@     �A@      K@      @      @      ;@      9@      @      @      A@      0@      &@      B@      9@     �D@      @      �?      �?      @      @      �?      @      @      �?      &@      &@      7@              @      :@      6@      @      @      =@      "@      $@      9@      ,@      2@      @              @      @      �?              1@       @      0@      �?      $@      *@                              �?      �?              �?       @      &@      �?      @      @                      @      @                      0@              @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��HThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?JZ��B@�	           ��@       	                    �?�2i�k+	@           h�@                          �<@:ވH}h@<           p~@                            @`0U��@           �z@������������������������       �D�m�|@�            0p@������������������������       ��I8x��@o            @e@                          �=@���)�>@!             M@������������������������       ����l�@             7@������������������������       �Z�%9�@            �A@
                           �?����w�	@�           ̑@                           �?[�Q� �@	            {@������������������������       ����-a@q            �f@������������������������       �O@		@�            `o@                           �?��|v��	@�           �@������������������������       ��TX#2	@�            �m@������������������������       �yG�:�	@6           `}@                            �?�Iq{�@�           ޡ@                          �3@Z9�qg~@p           ��@                           �?�8T蝣�?�             q@������������������������       ��i�c~ @H            �^@������������������������       �h1{By[�?Z            �b@                           �?�~���
@�            �r@������������������������       ��lc��j@6            �S@������������������������       ���'qX@�            �k@                          �4@s�h��S@G           ̚@                           �?��0�iG@;           ȋ@������������������������       ������� @�             s@������������������������       ��8�<@t           8�@                          �7@�mQ���@           Љ@������������������������       �]�2�@�            0x@������������������������       ���U��@           p{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     @r@     ��@      ?@      I@     0|@     �W@     @�@     `l@     X�@     @u@      @@      0@     `e@     �l@      4@      <@     �o@     �L@     �n@     @a@     �o@     `h@      3@       @     �M@     �P@      @      @      P@       @     �Z@      <@      X@     �G@       @       @     �K@     �L@      @       @     �H@       @     �Z@      9@     @V@      ?@       @       @      ;@      <@      �?              B@      @      Q@      1@      M@      0@       @              <@      =@       @       @      *@      @      C@       @      ?@      .@                      @      $@              @      .@                      @      @      0@                      @       @                      @                      �?       @      $@                               @              @      &@                       @      @      @              ,@      \@     @d@      1@      7@     �g@     �H@     `a@     �[@     �c@     �b@      1@      @      >@      P@      @      $@     @R@      0@     @S@     �@@     �N@     �K@      @       @      $@      ;@       @      @      I@      @     �A@      *@      *@      5@      �?      �?      4@     �B@      �?      @      7@      (@      E@      4@      H@      A@      @      &@     �T@     �X@      ,@      *@     �]@     �@@      O@     @S@      X@     @W@      $@      @      ?@      F@      "@              =@      (@      3@      9@      7@     �C@       @      @     �I@      K@      @      *@     @V@      5@     �E@      J@     @R@      K@       @      �?     @^@     �r@      &@      6@     �h@     �B@     ؈@     @V@     p�@      b@      *@              ?@     @P@       @      @      @@      *@     �l@      *@     @b@     �B@      �?               @      :@              �?      @             �`@      @     �T@      $@                       @      $@              �?      @             �L@      @     �B@      @                      @      0@                                     @S@      �?      G@      @                      7@     �C@       @       @      :@      *@     �W@      "@     �O@      ;@      �?                      ,@      �?      �?      $@      @      A@              (@       @                      7@      9@      �?      �?      0@       @     �N@      "@     �I@      9@      �?      �?     �V@     @m@      "@      3@     �d@      8@     ��@      S@     �y@      [@      (@             �D@      ^@      @      0@     �L@       @     0v@      7@     �k@     �H@                      0@      :@              @      .@             `d@      @     @P@      "@                      9@     �W@      @      "@      E@       @      h@      2@     �c@      D@              �?     �H@     �\@      @      @     �Z@      6@     `j@     �J@     �g@     �M@      (@              5@     �O@      �?       @     �H@      1@     �^@      @     �R@      5@      "@      �?      <@     �I@      @      �?      M@      @      V@      G@     @]@      C@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJzT�:hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��1��G@�	           ��@       	                   �8@�x�x �@�           ,�@                           �?�5hOV@�           �@                          �1@�Ҫoޚ@I           �@������������������������       ����@E            @Z@������������������������       ���t+�@            y@                          �2@D>�n�	@�           ,�@������������������������       �2�P�¹@�            �s@������������������������       ���#N�	@�           `�@
                           �?�A$�2�	@�           ��@                          �?@���V��@n            �f@������������������������       �/�m5��@e            �d@������������������������       ���qa@	             .@                          �;@E	��	
@4           �}@������������������������       �~��	g�	@�            `j@������������������������       ���ז�	@�            �p@                            �?E�ΐy�@-           ̚@                          �5@^�^j�"@�            �v@                          �1@Bk既� @�            @l@������������������������       ��I����?.             R@������������������������       ���3�9@e            @c@                           @�.>>E@T            �`@������������������������       ��t�R�}@7            @W@������������������������       ���:�@            �D@                          �6@��ȥ��@F           ,�@                           @�Z��P�@Z           `�@������������������������       �A��**@�            �i@������������������������       ��i���@�           ��@                           @�@9���@�            �w@������������������������       ���� @�             m@������������������������       ��F^7�f@W            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     ��@      =@     �J@     z@     @S@     ��@     �j@     ��@     0v@     �E@      3@     �k@     �u@      7@     �B@     �q@     �K@      w@     �e@     x@     �n@      A@      $@      b@     @p@      (@      9@      g@      A@     0s@     �W@     @s@      b@      .@             �H@     �R@               @     �E@      �?     @a@      2@     @a@     �D@                      @      2@                      (@             �E@      @      3@      @                     �F@     �L@               @      ?@      �?     �W@      ,@     �]@      B@              $@     �W@      g@      (@      7@     �a@     �@@      e@     @S@     @e@      Z@      .@      @      <@     �J@      �?       @      D@       @     �S@      7@      L@      @@              @     �P@     �`@      &@      5@     �Y@      ?@     �V@      K@     �\@      R@      .@      "@     �S@     �V@      &@      (@     @X@      5@     �O@     �S@     @S@      Y@      3@      �?      1@      =@       @      �?      :@       @      4@      3@     �A@      6@      @      �?      &@      <@              �?      9@      �?      4@      0@      A@      6@      @              @      �?       @              �?      �?              @      �?                       @      O@      O@      "@      &@     �Q@      3@     �E@      N@      E@     �S@      *@              @@      8@      @      @      =@      "@      =@      ?@      .@      9@       @       @      >@      C@      @      @      E@      $@      ,@      =@      ;@     �J@      @             @S@     �j@      @      0@     �`@      6@     h�@     �D@     {@     �[@      "@              2@      J@      @              ?@      @     @a@      $@      R@      >@                      @     �@@                      4@             �Z@      @      G@      ,@                              @                      @             �I@      �?      @      @                      @      ;@                      ,@              L@       @     �D@      &@                      .@      3@      @              &@      @      ?@      @      :@      0@                      @      .@      �?              &@      @      9@      @      0@      &@                      $@      @       @                              @      @      $@      @                     �M@      d@      @      0@      Z@      0@     �@      ?@     �v@      T@      "@              B@     @\@      @      "@     �P@       @     `z@      ,@     @o@     �E@      @              ,@      =@                      0@       @     @U@      @      F@      @      �?              6@      U@      @      "@     �I@             u@      $@     �i@     �C@      @              7@      H@              @     �B@       @     @W@      1@     �[@     �B@       @              2@      9@              �?      ;@      @      O@      @     �Q@      .@       @              @      7@              @      $@      @      ?@      $@      D@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?~���$H@�	           ��@       	                    �?��o~��@/           4�@                           �?wF`��p@�           ��@                           �?���q&�@�            �g@������������������������       ��F�m@.            �O@������������������������       ��n��o@V            @_@                          �6@��g$�@           �{@������������������������       ��wy� @�            @t@������������������������       �$�z�@E            �]@
                           @��#�@�           \�@                           @z�^*	@C           p@������������������������       �:YW���@           �{@������������������������       ����@&             M@                            @���Z@W            �@������������������������       �^pB-�@(           P}@������������������������       ����4� @/            �R@                           @�R��Ny@{           x�@                            �?�~cw��@Y           ��@                           �?UBn"�@�            @y@������������������������       �T��P�@@            @[@������������������������       � �<;V	@�            pr@                          �4@|X�t�@f           Ў@������������������������       �獦�6S@           �y@������������������������       ��_g	@_           ��@                          �7@uJ���@"           p�@                           @����M9@�           ��@������������������������       �R�����@q           ��@������������������������       �ۂFy@$            �I@                          �<@�h�~�@�            �k@������������������������       �8S唒�@h            �d@������������������������       �k/g�@%            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �s@     x�@      @@     �L@     0@      Q@     ��@      j@     ��@     �u@      :@      "@     �\@     �n@      1@      6@     �j@      4@     p|@     �S@     u@     �b@      ,@       @     �A@     @T@      @      @      H@       @     �o@      7@      `@     �D@       @       @      2@      =@      @       @      0@      �?     �F@      1@      ?@      6@       @       @      @      "@                      @              7@      @      *@      @                      ,@      4@      @       @      $@      �?      6@      ,@      2@      3@       @              1@      J@              @      @@      @      j@      @     @X@      3@                      @      C@              @      7@      @      e@      @      O@      ,@                      *@      ,@                      "@             �C@      @     �A@      @              @      T@     �d@      ,@      0@     �d@      (@     @i@      L@      j@     @[@      (@      @     �E@      V@      $@      @     �W@      $@     �K@     �H@     �P@     @P@      &@      @     �B@     �T@      "@      @     �S@      $@      K@     �A@      P@      L@       @              @      @      �?              0@              �?      ,@       @      "@      @       @     �B@     @S@      @      $@     �Q@       @     `b@      @     �a@      F@      �?       @     �B@     �P@      @      "@     �M@       @     �_@      @     �\@      D@      �?                      $@              �?      &@              4@              =@      @              .@     �h@     �q@      .@     �A@     �q@      H@     ��@      `@     `~@     �h@      (@      .@     �c@     �d@      *@     �@@     `k@      C@     �m@      [@      p@      a@      $@      @      F@      D@      �?      (@     �F@      1@      R@      B@     �T@      I@       @              0@      &@                      @              <@       @     �D@      @      �?      @      <@      =@      �?      (@      C@      1@      F@      A@     �D@     �G@      �?      (@     �\@     �_@      (@      5@     �e@      5@     �d@      R@     �e@     �U@       @      �?      >@     �C@      @      *@      R@       @     @W@      7@      X@      ?@       @      &@      U@     �U@       @       @     �Y@      *@     @R@     �H@     �S@     �K@      @              D@     �\@       @       @     �P@      $@     pr@      5@     �l@      O@       @              <@     @X@       @              =@      @      o@      @     �e@     �@@       @              ;@     �U@      �?              =@      @     �l@      @     `d@      :@                      �?      $@      �?                              2@       @      $@      @       @              (@      2@               @      C@      @      G@      ,@     �L@      =@                      &@      (@              �?      3@      @      D@      (@      H@      2@                      �?      @              �?      3@              @       @      "@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJR�*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?���p�0@�	           ��@       	                    @YF�Bf�@V           X�@                          �2@�X��)�@            �@                           �?E��D�@q             e@������������������������       �|>#-�@'            @P@������������������������       ��?���A@J             Z@                          �<@�d���8	@�           ��@������������������������       ��[��,	@m            �@������������������������       �������@>            �U@
                           �?�rW�@:           ��@                          �8@Ե��?�            �v@������������������������       �G��^i�?�             t@������������������������       �?A��@            �C@                          �1@r: g@b           h�@������������������������       ��}��/�@?            �X@������������������������       ����λ@#           �~@                           @���#Y@C           f�@                          �;@����.�@G           d�@                          �1@�yԡF#@�           ��@������������������������       ��pcw&s@e            �d@������������������������       ���x�ly@s            �@                           �?#�[U	@o             f@������������������������       ��9]e��@]            @b@������������������������       �ut�h�@             >@                           @����@�           Ј@                            @�����M@�           0�@������������������������       ���3�@�           �@������������������������       ��1g @O            �`@������������������������       �;z�0��@             4@�t�b��      h�h5h8K ��h:��R�(KKKK��h��B�
        4@     �q@     ��@      >@      N@     �|@     �R@     ȏ@     `l@     �@     �v@      3@      @      a@     @p@      0@     �A@     �k@      7@     �@     �X@     �t@      e@      @      @     @S@     @b@      (@      9@      ^@      5@     �b@      T@     �\@      [@      @       @      @     �@@       @              =@             �K@      @      7@      ,@              �?      �?      $@                      @              <@              &@       @              �?      @      7@       @              7@              ;@      @      (@      @               @      R@     @\@      $@      9@     �V@      5@      X@     �R@      W@     �W@      @             �P@     @W@      $@      6@     @T@      .@      W@     �O@     �U@     �R@      @       @      @      4@              @      $@      @      @      &@      @      4@              �?      N@     �\@      @      $@     �Y@       @     pv@      3@     @k@     �N@                       @     �E@                      5@      �?     �g@      @     �S@      *@                       @      @@                      4@              f@       @      R@      &@                              &@                      �?      �?      *@      @      @       @              �?      J@     �Q@      @      $@     @T@      �?      e@      *@     `a@      H@                      @      *@              @      @             �G@      @      5@      @              �?     �H@      M@      @      @      S@      �?     �^@      $@     �]@     �F@              .@      b@     �r@      ,@      9@     �m@     �I@     �@      `@     @}@      h@      ,@      .@     @Z@     @i@       @      8@      h@     �B@     `j@     �Z@      o@     �a@      (@      $@     �V@     @f@      @      ,@     @e@      =@     �h@      W@      m@     �X@      (@              0@      5@                      3@             �J@       @      B@      (@              $@     �R@     �c@      @      ,@     �b@      =@      b@      U@     �h@     �U@      (@      @      .@      8@       @      $@      7@       @      *@      ,@      1@     �F@              @      *@      ,@       @      @      3@       @      $@      $@      ,@     �F@                       @      $@              @      @              @      @      @                              D@     �X@      @      �?      G@      ,@     �r@      6@     `k@      I@       @              A@     �W@      @      �?      F@      (@     `r@      6@     @k@     �H@       @              >@      W@      @             �A@      &@     �m@      3@     �e@      D@       @              @       @              �?      "@      �?      M@      @      G@      "@                      @      @       @               @       @       @              �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJϢphG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @(���_@�	           ��@       	                   �8@_����@�           ¡@                          �3@��	?=@�           ��@                           @�LK@�           ��@������������������������       ������G@S           @�@������������������������       ���sR%�@i            `e@                           �?l~��+s@?           ��@������������������������       ���М@�            �m@������������������������       �<^�{�@�           P�@
                           �?ܻ �	@�           ��@                           @�ߝ���	@P           �@������������������������       ��v̅	@.           �|@������������������������       ��b�ՏO@"             K@                           �?>6 �y�@T             ^@������������������������       �����@             A@������������������������       �W���@�@>            �U@                           @k��=h@2           ��@                          �4@���@�            �w@                           �?v�7��@�            @i@������������������������       �
��@J            @\@������������������������       �uv?'8�@=            @V@                           �?UU���@r            �e@������������������������       �qB~f�P@;            �X@������������������������       �Q|�g@7            @S@                           �?'sK3��@9           ��@                            @�E?� @           �{@������������������������       ���°��@�            0v@������������������������       �?�]Κ�?4             W@                            �?n �Wq�@           ��@������������������������       ��i6v�@v            �f@������������������������       �켿#@�           ؃@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     @�@      6@      H@     �{@     �W@     p�@     �l@     �@     x@      >@      0@     �j@     �t@      2@      B@     s@     �Q@     �x@      h@      y@     �p@      9@      "@     `b@     �m@      (@      6@     �l@     �A@     pt@     @\@      t@     �e@      0@      @      G@     �W@      @      @      S@      (@     `f@     �I@     @c@     �V@      @      @      >@      K@      @      @     �K@      "@     �b@      A@     �`@     @S@              �?      0@     �D@      �?              5@      @      >@      1@      6@      ,@      @      @     @Y@      b@       @      0@      c@      7@     �b@      O@     �d@     �T@      &@              <@     �A@      @      �?      <@      �?     �O@      $@     �K@      *@              @     @R@     @[@      @      .@      _@      6@     @U@      J@     �[@     �Q@      &@      @     @P@     �W@      @      ,@     @S@     �A@     �P@     �S@      T@     @X@      "@      @     �H@     �R@      @      (@     @Q@      ;@     �I@      P@     �N@      U@      @      @      G@     @Q@      @      (@     �O@      6@     �C@      I@     �N@     �S@      @       @      @      @      �?              @      @      (@      ,@              @      �?              0@      5@               @       @       @      0@      .@      3@      *@       @              @      @                              @      @      @      @      @       @              (@      2@               @       @      @      "@      &@      (@      $@                     �Y@     @k@      @      (@     `a@      9@      �@      C@      y@     �\@      @              >@      O@               @      9@      1@     �^@      "@      S@      <@      @              7@     �C@                       @      @     �R@      @     �C@      &@                      ,@      2@                      @             �D@      @      3@      $@                      "@      5@                       @      @     �@@              4@      �?                      @      7@               @      1@      ,@     �H@      @     �B@      1@      @               @      @               @      (@      &@      <@              1@      .@      @              @      1@                      @      @      5@      @      4@       @                     @R@     �c@      @      $@     �\@       @     �|@      =@     `t@     �U@                      &@     �L@                      :@       @     �j@      $@     �[@      3@                      "@      L@                      6@       @     �c@      "@     �T@      0@                       @      �?                      @             �J@      �?      <@      @                      O@     �X@      @      $@      V@      @     �n@      3@      k@     �P@                      4@      2@              �?      .@      @     @Q@      @      E@      "@                      E@     @T@      @      "@     @R@      @      f@      .@     �e@      M@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��?$(w@�	           ��@       	                    �?������@z           Z�@                           �?����č@�           �@                            �?�0�-"@:           ~@������������������������       ���_��@`             a@������������������������       �y��ӹ?@�            �u@                            �?jq��@p             h@������������������������       ������r@E            @]@������������������������       ���}>�@+            �R@
                           �?nUa��	@�           0�@                           �?9�ZW�	@�           ��@������������������������       ���	}@�            �x@������������������������       � �j�
@�           ��@                          �5@+o9��@           �y@������������������������       ��`��vN@�            `l@������������������������       ����@y            �g@                          �4@<��_�,@+           p�@                           �?�R��G6@B           (�@                            @�E�n�]@@           �@������������������������       ��Ey��%@           0{@������������������������       �VE{�;�@/            �R@                           @0�>]��@           pz@������������������������       ���S��?�            Ps@������������������������       ��C�@E            �\@                           @7eC<_�@�           ��@                          �8@��fo�@X           �@������������������������       �u��U0@�            s@������������������������       �Lw;��@�            �i@                          �9@$�$�%@@�             o@������������������������       �M���%@f            �e@������������������������       ���H�	U@+            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �q@     ؀@      >@      N@     p~@     �S@     8�@     �k@     ��@      w@      A@      7@     �h@     �s@      4@     �H@     �u@      P@     v@     �f@     y@     @n@      <@       @      M@     �T@      �?      $@      T@      $@     �d@      D@     `d@     �M@      �?       @      G@      R@      �?      "@      N@      @     �X@      @@     @Z@      I@      �?       @      ,@      8@                      2@       @      :@      @     �B@      "@                      @@      H@      �?      "@      E@       @     @R@      ;@      Q@     �D@      �?              (@      &@              �?      4@      @     �P@       @      M@      "@                       @      @              �?      @       @     �G@       @     �D@      @                      @      @                      *@      @      4@      @      1@      @              5@     �a@     �l@      3@     �C@     �p@      K@     `g@     �a@     �m@     �f@      ;@      5@     �[@     �d@      3@      8@     @j@      C@     �\@     �Z@     �c@     �a@      :@      @      3@     �R@      @      *@     �S@      @      I@      ?@      N@     �J@      @      0@     �V@      W@      ,@      &@     �`@      @@      P@      S@     �X@     �U@      6@              >@     �O@              .@     �M@      0@     @R@     �A@      T@     �E@      �?              @      B@              (@      9@      @      O@      3@     �G@      0@                      8@      ;@              @      A@      (@      &@      0@     �@@      ;@      �?             �U@     `l@      $@      &@     @a@      .@     0�@      D@      z@      `@      @              C@     @`@      @      @     �H@      @      y@      .@     �l@     �M@                      5@      O@      @      @     �C@             �l@      @     @[@     �B@                      4@      M@       @      �?      >@              i@      @     �T@      A@                      �?      @       @       @      "@              <@              :@      @                      1@      Q@              �?      $@      @     �e@       @     �]@      6@                      *@      L@              �?      @      @     ``@             @W@      @                      @      (@                      @             �E@       @      :@      1@                     �H@     @X@      @      @     @V@      &@     �j@      9@     �g@     @Q@      @              4@      R@      @      @     �L@      "@      d@      *@     ``@     �C@                      ,@     �G@      @              A@       @     �Y@      @     �R@      2@                      @      9@              @      7@      �?     �L@      "@     �L@      5@                      =@      9@      @      �?      @@       @      J@      (@     �L@      >@      @              3@      7@      @              ,@      �?     �F@      "@      ?@      7@      @              $@       @              �?      2@      �?      @      @      :@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�2dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����)u@�	           ��@       	                    �?��^5��@l           :�@                          �2@��ԣ?Q	@           ԙ@                           @4��t��@�            �s@������������������������       ����OF�@�            �o@������������������������       ���� �@*             P@                          �4@�W%�:�	@8           ܔ@������������������������       ��Õ(�a	@�            �r@������������������������       ��J�n�	@�           $�@
                           �?�&�tA@h           @�@                            �?��d
�@�             k@������������������������       ������@*            �O@������������������������       ���z��@c             c@                            �?,���*x@�             u@������������������������       ����<�@|            �f@������������������������       �ȁ��F@_            @c@                          �7@ޘd@=           ��@                           @��=n@?           ��@                           �?�<n�|�@�            �t@������������������������       �G�%b+�@h            @e@������������������������       ��{���� @]            `d@                           �?��Ex|@z           ��@������������������������       ��6/ԣ��?�            �t@������������������������       �r���@�            �@                           @�rT*��@�            �x@                           �?��{:�@�            Pu@������������������������       �t��G)@C             [@������������������������       ��5K�@�             m@                           @���g��@#            �K@������������������������       ��#�Z�n@             6@������������������������       ��ND��F@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      q@     �@     �C@     �K@     �~@     �T@     ؎@      l@     ��@      x@      ;@      2@      i@      u@      =@      E@     �t@     �N@      v@     �f@     �u@     �q@      9@      2@     �c@      o@      =@     �@@     �o@     �G@     �m@     @`@     �n@     �l@      8@      @      9@      E@      �?       @     �K@              Q@      8@      L@     �D@               @      .@      <@      �?      �?     �H@             @P@      0@     �I@      :@               @      $@      ,@              �?      @              @       @      @      .@              ,@     �`@     �i@      <@      ?@     �h@     �G@      e@     �Z@     �g@     �g@      8@       @      :@      =@       @       @     �F@      (@      I@      2@     �G@      I@      *@      (@     �Z@      f@      4@      =@     @c@     �A@     �]@      V@     �a@     `a@      &@              E@      V@              "@     �R@      ,@     �]@      I@     �Y@      J@      �?              $@     �A@              �?     �@@      @     �D@      6@     �F@      8@                       @      .@                      ,@      �?      *@      @      &@      @                       @      4@              �?      3@      @      <@      2@      A@      5@                      @@     �J@               @      E@      "@     @S@      <@      M@      <@      �?              4@      9@              @      .@      @     �F@      *@     �E@      $@      �?              (@      <@              @      ;@      @      @@      .@      .@      2@              �?     �R@     @n@      $@      *@      d@      5@     ȃ@      F@     @y@      Z@       @             �I@     `h@      "@      @      Y@      ,@     �@      6@     s@     �P@      �?              3@     �L@       @              6@      (@     ``@       @     @P@      1@                      ,@      ?@                      0@      $@     �I@      @      >@      &@                      @      :@       @              @       @      T@      �?     �A@      @                      @@     @a@      @      @     �S@       @     �y@      ,@      n@      I@      �?              "@     �D@      �?              1@              g@      @     @Q@       @      �?              7@     @X@      @      @     �N@       @      l@      $@     `e@      E@              �?      7@     �G@      �?      @      N@      @      W@      6@     �X@     �B@      �?      �?      (@      C@              @     �I@      @      U@      1@     @W@      A@                      �?      *@                      &@      @      :@      @      E@      @              �?      &@      9@              @      D@              M@      ,@     �I@      ;@                      &@      "@      �?              "@       @       @      @      @      @      �?              �?      @                      @              @              @      @      �?              $@      @      �?              @       @      �?      @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�{eBO�@�	           ��@       	                    �?�"��	@�           Ę@                           �?������@)           @}@                          �4@�I���@�            �k@������������������������       �'-fo��@;            @V@������������������������       �\���@R            ``@                            �?2�NB��@�             o@������������������������       �n���p @2            @R@������������������������       �  ���@j            �e@
                          �:@_��o��	@�           t�@                           @~陇�]	@/           ��@������������������������       �pXdL�[@`           ��@������������������������       �&��َ�	@�            ps@                          @@@�
F	@�            �p@������������������������       �TdP��	@�            @l@������������������������       �}�ɔ�V@             C@                          �4@�+B�@�           0�@                           @�� (��@�           Ē@                          �2@������@�            �q@������������������������       �L4�P�@c            �b@������������������������       ��Zg�%�@S            �`@                           �?�_��@A           ��@������������������������       �B��3�?�            �t@������������������������       �ݱ0C@o           8�@                           @8���@�           ��@                           @\�}@�@�           ��@������������������������       �ZնV�@2           �~@������������������������       �@�ɐk@x           ��@                          �:@Y�I�@             D@������������������������       �*�9	�@             <@������������������������       �η:�?             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `p@     0�@      =@     �G@     �{@      T@     x�@     �h@     0�@     �v@      ?@      1@     �a@     �l@      0@      >@     `m@     �F@     �m@     �]@     �q@     `i@      :@       @     �C@     �Q@       @       @      Q@       @      Z@      4@      [@      E@       @       @      4@     �C@       @      @     �A@       @     �H@      (@     �A@      0@      �?              @      ,@                      &@      �?     �@@      @      (@      "@      �?       @      1@      9@       @      @      8@      �?      0@      @      7@      @                      3@      @@              �?     �@@             �K@       @     @R@      :@      �?              @      0@                      $@              @              ?@      @      �?              .@      0@              �?      7@              H@       @      E@      6@              .@     �Y@      d@      ,@      6@     �d@     �E@     �`@     �X@     �e@      d@      8@      "@     �R@     �a@      &@      3@     ``@      ;@     @]@      R@      a@     �X@      1@       @     �E@     �Q@      @      $@     @W@      5@     @V@      =@      Z@     �Q@      @      @      @@     �Q@      @      "@      C@      @      <@     �E@     �@@      ;@      *@      @      <@      4@      @      @      B@      0@      1@      ;@      C@     �O@      @      @      6@      0@      @      @      A@      0@      *@      7@      A@     �H@      @              @      @                       @              @      @      @      ,@              �?      ^@     �s@      *@      1@      j@     �A@     ��@      T@     X�@     �c@      @              F@     �c@      @      &@      R@      @     �@     �B@     `r@     @P@       @              .@     �@@      @      @      <@             @V@      3@     �R@      2@                      @      0@              �?      0@             �L@      $@      A@      &@                      $@      1@      @       @      (@              @@      "@     �D@      @                      =@      _@      @       @      F@      @      z@      2@     `k@     �G@       @              $@      C@               @      "@             @g@      @     @S@      @       @              3@     �U@      @      @     �A@      @      m@      ,@     �a@      D@              �?      S@     @d@      @      @      a@      >@     Ps@     �E@     Pp@     @W@      @      �?     �P@      d@      @      @     @`@      :@     0s@     �A@      p@     �V@      @      �?     �E@      Q@              @      Q@      4@     @]@      2@      Z@      F@      @              7@      W@      @      @      O@      @     �g@      1@     @c@     �G@                      $@       @       @              @      @       @       @      @       @                       @       @       @              @      @       @       @      @       @                       @                              @      �?                                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ۺKhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �7@��q�o@�	           ��@       	                    �?��=(:@�           H�@                            @妣8U�@�           �@                           @o�sS@&           ��@������������������������       �3e�abi@!            }@������������������������       ��jy�g�@            z@                          �2@��Z95�@�            �t@������������������������       �0O���L@P            @a@������������������������       ����N�@w            �g@
                           �?�O���@�           ��@                          �2@�h�B�>@           P{@������������������������       ��A͙��@u            �f@������������������������       �V9[�{@�            �o@                           @?�ֻr�@�           А@������������������������       �f����@�           h�@������������������������       ����L��@�            pz@                          �;@�5*�@	@�           ��@                           @ܶ�$܇@�           ��@                          �:@O
Ɋ�	@$           �|@������������������������       �_	v�wO	@�            �v@������������������������       ��W+��@9            @W@                          �8@�	ڌ@�            �p@������������������������       �ƳQq+z@A             Y@������������������������       ������@p            �d@                           @ݑ��Z{	@           }@                           �?l���	@�            0t@������������������������       ���@2             Q@������������������������       �n\EcGq	@�            �o@                            @^;Lu)W@T            �a@������������������������       �4�+�r@C            �[@������������������������       �|e�3�G@             ?@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �r@     ��@      C@      M@     �{@     �Q@     ��@     `j@     ��@     �x@      >@      $@     �g@     0z@      1@     �B@     �r@      A@      �@     @Z@     @�@     �j@      .@       @     �T@     �i@      "@      $@      b@      *@     �w@      @@      m@     �X@      @      �?      M@     �a@      @      @     @[@      *@     @r@      :@     �d@      N@      @      �?      C@     @V@       @      @     �M@      *@     @[@      8@     @S@      F@      @              4@      K@      �?              I@             �f@       @     �V@      0@              �?      8@     �N@      @      @      B@              V@      @     @P@      C@                       @      8@       @              (@              I@      �?      ?@      $@              �?      0@     �B@      @      @      8@              C@      @      A@      <@               @     @[@     �j@       @      ;@      c@      5@     @z@     @R@      v@     @]@      &@             �C@     �Q@      �?              >@             `b@      &@     �]@      2@      �?              @      6@                      (@              U@      @      E@       @      �?              @@     �H@      �?              2@             �O@      @     @S@      $@               @     �Q@      b@      @      ;@     �^@      5@     q@      O@      m@     �X@      $@       @     �G@     �U@      @      7@     �V@      0@      ]@      L@     �_@     �Q@      "@              7@      M@       @      @      @@      @     �c@      @     �Z@      =@      �?      .@     @Z@     �b@      5@      5@      b@      B@     �g@     �Z@     �i@     �f@      .@      @     �N@      W@      "@      (@     @W@      *@     �b@     @Q@     �`@     �S@      (@              E@     �Q@      "@      @      Q@      *@     �P@      J@      P@      L@      (@             �@@      O@       @      @     �J@      *@     �G@     �D@      K@     �B@      &@              "@       @      �?              .@              3@      &@      $@      3@      �?      @      3@      6@              @      9@             �T@      1@     @Q@      6@              @      @      "@                      0@              ;@      @      9@      @                      (@      *@              @      "@             �K@      (@      F@      .@              &@      F@      L@      (@      "@      J@      7@     �E@     �B@      R@     �Y@      @      &@     �@@     �@@      (@       @      <@      6@      0@      =@     �G@     @T@      @       @      @       @      @      �?      $@              "@      @      (@      ,@              "@      >@      9@      "@      @      2@      6@      @      7@     �A@     �P@      @              &@      7@              �?      8@      �?      ;@       @      9@      6@                      $@      5@                      3@      �?      .@      @      6@      1@                      �?       @              �?      @              (@       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJୋ_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @ra�Wk@�	           ��@       	                    �?{�GA�@}           ��@                           �?_���@�           �@                          �<@���$>�@,           @~@������������������������       �5z���@           `z@������������������������       ���SO��@(             O@                           �?)��ǖG@t            �g@������������������������       ���,YH�@7            �V@������������������������       �4�i��@=            @Y@
                          �3@��L�|	@�           И@                           @~���Ŷ@,           �}@������������������������       �//�E@d@!           �|@������������������������       ����RǸ@             .@                           @ٿk�e�	@�           l�@������������������������       ���DN�	@R           ��@������������������������       ��?p�@_            �c@                           �?%z52�@%           ș@                           @�{r�� @h           X�@                            �?R)=gr��?�            �v@������������������������       ���;��?9            @U@������������������������       ����4C�?�            pq@                          �4@x/����@|            �g@������������������������       �z�;���@?            @W@������������������������       ��[�3u}@=            �X@                           @�=P��x@�           �@                          �4@����8@�            �@������������������������       ��=��1�@           �x@������������������������       �4�M+K�@�            @w@                           @�x�)L�@�            pt@������������������������       �<���fa@(             Q@������������������������       �M��Le[@�            0p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �r@     ��@      D@     �Q@     �}@     �Q@     Ȏ@      l@      �@     w@      =@      &@     �l@     @u@      ?@      H@     t@     �J@     `v@     �g@     �y@      o@      :@              Q@      X@       @      "@     @U@      @      d@      @@      d@      M@      �?             �I@     @S@       @      "@     �P@      �?      Y@      >@     �X@     �H@                     �G@      R@       @      @     �K@      �?     �X@      7@     �V@      >@                      @      @              @      &@              �?      @      "@      3@                      1@      3@                      3@       @     �N@       @     �N@      "@      �?              @      ,@                      $@      �?     �@@              5@      @                      $@      @                      "@      �?      <@       @      D@      @      �?      &@     @d@     �n@      =@     �C@     �m@      I@     �h@     �c@      o@     �g@      9@      @     �B@      N@              @     �P@      &@     @X@     �I@     �V@      I@      @      �?     �B@     �M@              @      O@      $@     �W@     �I@      V@     �H@       @       @              �?                      @      �?       @               @      �?       @       @     @_@      g@      =@     �A@     @e@     �C@      Y@     @Z@     �c@     �a@      5@      @     @Z@     �b@      <@      >@      c@     �B@      U@     @T@     �b@      ^@      1@      @      4@      B@      �?      @      2@       @      0@      8@       @      5@      @      �?     @R@     �g@      "@      6@     �c@      1@     ��@      B@     �x@      ^@      @              (@      R@               @     �C@      �?     pp@      @     �a@      5@      �?              @      D@                      7@      �?     �h@       @      V@      $@                              *@                      @      �?      K@              (@       @                      @      ;@                      4@             �a@       @      S@       @                       @      @@               @      0@             �P@      �?     �J@      &@      �?               @      &@               @      @             �C@              6@      @      �?                      5@                      &@              <@      �?      ?@      @              �?     �N@     �]@      "@      4@     @]@      0@     �v@     �@@     �o@     �X@       @      �?     �D@     �U@       @      @      T@      @     �q@      ,@     �e@      R@      �?              *@      H@              @      4@       @     �c@       @      X@     �G@              �?      <@     �C@       @      @      N@      @      _@      @     �S@      9@      �?              4@      ?@      @      *@     �B@      $@     �T@      3@      T@      ;@      �?               @      @       @       @       @      @      ,@      &@      @      &@                      2@      ;@      @      &@      =@      @      Q@       @     @R@      0@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��V[Y@�	           ��@       	                    @Vu�Jq�@h           *�@                           �?В|�c�@�           |�@                            �?����}@�            @v@������������������������       ��gnL�@E            �]@������������������������       ��&C/;�@�            �m@                           �?Y6w�~@�           ؇@������������������������       �����@�            �q@������������������������       ����8^@1           �}@
                           @���o2@�           ؐ@                           @W�^	��@�            `n@������������������������       ����'�@�             i@������������������������       ������@             E@                           @�����t@           �@������������������������       �<��") @R            �@������������������������       ��ӎ�`S@�            �q@                            �?s5F�%�@P           К@                           @|4�9�Q	@2           �}@                           �?�2�K��	@�            pt@������������������������       �ͭ�g�@7            @X@������������������������       ���	@�            �l@                           �?��HV�\@`             c@������������������������       �]e�m�8@+            �Q@������������������������       ���v���@5            @T@                           @
���"R@           T�@                          �:@D�@�           H�@������������������������       ��#j�*@>           @������������������������       �HA�E��@�            �q@                           @��az�@&           �|@������������������������       �N#	>@�            0p@������������������������       ���(�P@�             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     ps@     ��@      ?@      L@      {@      S@     ��@     @l@     �@     `x@      =@      @      ^@     �r@      ,@      6@     `i@     �B@     X�@     �Z@     ��@     �d@       @      @     �S@     �d@      $@      *@     �a@      :@      m@     @W@     �k@     �^@      @              ?@     �J@      �?      @     �B@      @     �X@      *@      V@      :@                      @      7@              �?       @       @      8@      @      F@      "@                      ;@      >@      �?      @      =@       @     �R@      "@      F@      1@              @      H@     @\@      "@      "@     �Z@      6@     �`@      T@     �`@      X@      @      @      1@      N@      @       @      B@      $@      H@      ?@      B@     �A@      �?      @      ?@     �J@       @      @     �Q@      (@     �U@     �H@     �X@     �N@      @             �D@     �`@      @      "@      N@      &@      |@      *@     @s@     �F@      @              2@      B@                      *@      "@     �S@      @      R@      &@      �?              .@      <@                      *@      "@     �P@              O@      @                      @       @                                      (@      @      $@      @      �?              7@     �X@      @      "@     �G@       @     0w@      "@     �m@      A@       @              1@      N@       @       @      6@             pp@      @     �c@      4@                      @      C@       @      @      9@       @      [@      @      T@      ,@       @      &@     �g@     �l@      1@      A@     �l@     �C@     �r@      ^@     �r@     �k@      5@             �H@     �L@      "@      1@     �N@      ,@      T@     �E@     @T@     �M@      "@             �B@      B@      @      1@      H@      *@     �D@      A@      H@      D@      "@              @      $@              @      .@              5@      0@      ,@      @      @              >@      :@      @      (@     �@@      *@      4@      2@      A@      A@      @              (@      5@      @              *@      �?     �C@      "@     �@@      3@                       @      ,@                      @              ,@      @      2@      @                      @      @      @               @      �?      9@      @      .@      *@              &@     �a@     �e@       @      1@     @e@      9@      k@     @S@     �k@     �d@      (@      $@     @^@     �\@      @      &@     �[@      3@     @U@     �O@     @[@     @]@      &@             �S@     �V@      @       @     @S@      (@      K@     �B@     @S@      K@       @      $@      E@      8@              "@     �@@      @      ?@      :@      @@     �O@      @      �?      5@      M@      �?      @      N@      @     �`@      ,@     @\@     �G@      �?      �?      @      ?@              @      2@      @      X@      "@     �O@      9@                      1@      ;@      �?              E@              B@      @      I@      6@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJq�bmhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�[[z��@�	           ��@       	                    �?�k��@|           l�@                          �1@L��i�@U           ��@                           �?P��M5�?�             n@������������������������       ��3�OW� @)             R@������������������������       �S��[�?r             e@                           @J�ֿ�@�            �r@������������������������       �-����@q            �f@������������������������       �W8k%�?I            �]@
                           @'2ٱ�@'           ��@                          �2@��EA@T           ��@������������������������       �(�%6�@�            `x@������������������������       ���*S�@e            �e@                          �1@��oS�q@�            �t@������������������������       ���ɷ�� @]             b@������������������������       ��ae��@v            @g@                          �;@}�5ٷ�@           \�@                           �?�s^8@           �@                           �?8����@q           �@������������������������       ���(@�            0u@������������������������       ���b��@�            �p@                           @��k��@�           ��@������������������������       ���p�w�@           ��@������������������������       �<�`�@w            �g@                           �?��c�C	@           �y@                          �=@Vj<X^	@�            �m@������������������������       �e����@P            @\@������������������������       �;^*�k@P            �_@                          �=@Z����Z@q             f@������������������������       �O#f�{@:            �V@������������������������       ���:@7            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      s@     H�@     �A@     �M@     p}@     �R@     ��@     @l@     `�@     �w@     �B@      @     �R@     �d@      @      (@     @]@      .@     8�@      K@     �u@     �^@      �?              <@     �K@              @     �@@       @      o@      @     �`@      @@                      $@      5@              �?      3@              `@              K@       @                       @      @                      &@             �A@              (@      @                       @      ,@              �?       @             @W@              E@      @                      2@      A@               @      ,@       @      ^@      @     @T@      8@                      .@      7@               @      ,@       @     �E@      @     �M@      4@                      @      &@                                     @S@       @      6@      @              @      G@     @[@      @      "@      U@      *@     �p@     �G@     �j@     �V@      �?      @      C@     �R@      @      @     �O@      *@     �b@      F@     �W@     @R@      �?      @      ;@      L@      �?             �I@      @     �X@      =@     �Q@      H@              �?      &@      2@       @      @      (@      @      I@      .@      9@      9@      �?               @     �A@      �?      @      5@             �^@      @     �]@      2@                      @      3@              @      @              L@      �?     �I@      @                      @      0@      �?              ,@             �P@       @     �P@      .@              ,@     �l@     Px@      ?@     �G@      v@      N@     �|@     �e@      {@     �o@      B@      @     `f@     �t@      :@      A@     �q@     �F@     {@     `a@      w@     �f@     �@@              J@     �X@      �?      @     �S@      @      g@      =@     @]@     �A@      @              :@     �J@              @     �G@      �?     @^@      0@      H@      2@       @              :@     �F@      �?              @@      @     �O@      *@     @Q@      1@       @      @     �_@     �m@      9@      ;@     �i@     �D@      o@     �[@     `o@     `b@      =@      @     @Z@     �h@      3@      ;@     �f@     �C@     @k@     @T@     �m@     �`@      7@       @      6@     �C@      @              8@       @      ?@      =@      ,@      ,@      @      "@     �I@     �K@      @      *@     @Q@      .@      9@     �@@      P@     @R@      @      "@      C@     �@@      @      $@      A@      *@      @      5@      8@     �G@       @      @      ,@      $@       @      @      &@      $@      @      @      .@      A@      �?      @      8@      7@      �?      @      7@      @       @      1@      "@      *@      �?              *@      6@       @      @     �A@       @      4@      (@      D@      :@      �?              @      2@                      ,@              *@      @      <@      "@                      "@      @       @      @      5@       @      @      @      (@      1@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�UPhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �1@=P�t@�	           ��@       	                    �?�ՄEA@p           ȁ@                           �?y�;�ku @�             m@                            �?Pq��v� @M             ^@������������������������       ���9Z� @+            �P@������������������������       ���v3_�?"             K@                            �?��k���?L             \@������������������������       �%��G�?             ;@������������������������       ��(�!<& @;            @U@
                           @󉔏i�@�            u@                            �?�R�V�%@h            �d@������������������������       ���>9�@4            �U@������������������������       ���Dd@4             T@                           @��d��X�?o            @e@������������������������       ���)Z�?J             [@������������������������       ��컪@�?%             O@                           �?����@>            �@                           �?��'�;�	@�           h�@                           �?�ό�@           �y@������������������������       ����M@`            �b@������������������������       ��4�b�B@�            �p@                            �?iw�h�F
@�           ��@������������������������       ��=Sv`M	@�            �r@������������������������       ��)pr�
@�           ��@                           �?�N@�2�@�           ؝@                           @���U@p           ��@������������������������       �u��u�@h            �e@������������������������       �<�	C��@           �z@                          �<@w����@?           x�@������������������������       �n�$풓@           ��@������������������������       ���e��@=             X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        =@     Ps@     ȁ@     �A@      M@     �z@      U@     ��@     �j@     0�@      t@     �C@       @      9@     �U@                      @@             @o@      5@     �]@     �@@                      $@      6@                      6@             @^@      @     �F@       @                      @      *@                      ,@             �O@       @      2@      @                      @      &@                      $@              @@              @       @                               @                      @              ?@       @      &@      @                      @      "@                       @              M@       @      ;@       @                              @                                      1@      �?      @                              @      @                       @             �D@      �?      7@       @               @      .@     @P@                      $@              `@      1@     �R@      9@               @      ,@      B@                      @             �G@      ,@      :@      6@               @      @      5@                                      3@      &@      *@      ,@                      @      .@                      @              <@      @      *@       @                      �?      =@                      @             �T@      @      H@      @                      �?      0@                      @             �H@             �A@      @                              *@                                     �@@      @      *@                      ;@     �q@      ~@     �A@      M@     �x@      U@      �@     @h@     x�@     r@     �C@      9@     `d@      h@      7@     �C@      l@      I@     �g@      ^@     �l@     `b@      <@      �?     �L@      N@      @      $@      C@      @      U@      3@     @V@     �E@      @      �?      4@      3@                      ,@             �D@      @      B@      (@      �?             �B@     �D@      @      $@      8@      @     �E@      .@     �J@      ?@       @      8@     �Z@     �`@      4@      =@     @g@     �F@     �Z@     @Y@     �a@      Z@      9@      @      B@     �B@       @      @      O@      "@      B@     �A@      F@      2@      $@      3@     �Q@      X@      2@      7@      _@      B@     �Q@     �P@     �X@     �U@      .@       @     @^@     r@      (@      3@      e@      A@     (�@     �R@     �|@     �a@      &@              ;@     �S@       @       @      A@      @     `p@      ,@     `b@      <@      �?              &@      4@               @      2@      �?     @Q@      @     �C@       @      �?              0@     �M@       @              0@      @      h@      $@      [@      4@               @     �W@     @j@      $@      1@     �`@      >@     �s@      N@     Ps@     �\@      $@       @     @S@     �h@      $@      .@     �\@      ;@     Ps@     �K@     �r@     �W@      $@              1@      (@               @      4@      @      $@      @       @      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��r`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�IN�]R@�	           ��@       	                    �?Z,�	@�           ��@                          �<@j����@�           P�@                           �?�DzI	>@X           Ѐ@������������������������       ���c��@p            �e@������������������������       ��@�            �v@                          �>@I��V�9@*             T@������������������������       �GQGɼ$@            �D@������������������������       ���^$�@            �C@
                           �?� ���	@f           ��@                          �1@�*���	@�             w@������������������������       ��N�w�!@             =@������������������������       ��o�>�	@�            Pu@                            �?�l!J.4	@�           �@������������������������       �[	o�Y@u             h@������������������������       �>a
�`	@            z@                          �4@K�Z�=C@�           �@                           @<��Ȼc@�           t�@                           @ �'X��@*           �|@������������������������       �U�6�Q@�            Pv@������������������������       �$=�P�@E             Y@                           @{ˣ{��@�           ��@������������������������       ��O0��� @7           �@������������������������       �#ǴP�@�            `k@                           �?�׫@�           ��@                          �=@2���Q@�             s@������������������������       ���)��M@�            �q@������������������������       �:z�0��@             4@                          �5@/'�ƫ@           �@������������������������       ��ǨW�@V            �`@������������������������       �XVS��@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     0s@     ��@      @@     �G@     �}@     @R@     H�@     �l@      �@     �v@     �A@      1@     �e@     @k@      1@      :@     �o@     �F@     �m@     �`@     p@     �h@      9@      @      I@     �U@       @      "@     @X@      @     ``@      B@      \@     @S@      "@      @      B@     �R@       @      @     �V@      @     �_@     �@@     �X@     �K@      "@      �?      &@      1@                      :@             �M@      @      G@      "@       @       @      9@     �L@       @      @     @P@      @     �P@      >@     �J@      G@      @              ,@      *@               @      @       @      @      @      *@      6@                      @      *@               @      @      �?      �?      �?      @      $@                      "@                              @      �?      @       @       @      (@              ,@     �^@     ``@      .@      1@     �c@      D@     @Z@     @X@      b@     �^@      0@      @     �D@     �M@      &@      @      H@      7@      H@      C@      C@     �I@      @      �?              @      @                              @      @      @      @               @     �D@     �K@       @      @      H@      7@     �F@     �@@      @@      F@      @      &@     @T@      R@      @      *@     @[@      1@     �L@     �M@     �Z@     �Q@      $@              >@      8@      �?      @      ?@       @      *@      3@     �C@      6@       @      &@     �I@      H@      @      "@     �S@      "@      F@      D@      Q@     �H@       @      �?     �`@     �s@      .@      5@     `k@      <@     �@      X@     ��@     `d@      $@             �K@      d@      @      &@     @T@      @     �}@     �E@     �p@     �Q@                      ;@     �R@       @      @      C@       @     `d@      ?@     �S@     �B@                      4@      I@       @      @      A@      �?     �a@      ,@     �N@      >@                      @      9@                      @      �?      6@      1@      1@      @                      <@     @U@      @      @     �E@      �?     �s@      (@      h@      A@                      7@     �J@              @      >@             �n@      (@      ^@      1@                      @      @@      @      @      *@      �?     @Q@             @R@      1@              �?      T@     �c@       @      $@     @a@      9@     �q@     �J@      q@      W@      $@              @      I@      �?              =@             �\@      @     @T@      *@      �?              @      I@      �?              5@              \@      @      T@      $@                                                       @              @      @      �?      @      �?      �?     @R@      [@      @      $@     @[@      9@     `e@      G@     �g@     �S@      "@              @      0@               @       @      "@      =@      @      G@      "@      @      �?     �Q@      W@      @       @     @Y@      0@     �a@     �D@      b@     �Q@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�� `hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?R2�.@�	           ��@       	                   �3@_��b;@           ��@                           @��u��j@\           �@                           �?+LХ�@�            �o@������������������������       �jq=�p@n            �e@������������������������       ���U�@0            @T@                           @�{����?�            `r@������������������������       �'�3)��?`            �b@������������������������       ��.ke�?^            �a@
                          �<@M��x�@�           ��@                           �?u���`@@�           ��@������������������������       ����;��@�            �p@������������������������       �����T@�            �v@                           @���+�D@2             R@������������������������       �-�{4S@$            �J@������������������������       ����bH @             3@                           @
�9z�(@�           Ф@                           �?�q��Vm	@�           \�@                           @<�ѺF�	@S           ��@������������������������       ��x�J҄@6            �V@������������������������       �.�N3Np	@           �{@                            �?gX/�(	@�           �@������������������������       ���ϮL	@_           �@������������������������       �u�9��@/            ~@                           @��{�'@�           D�@                            @���@�@�           ��@������������������������       �|�bh�-@�           Ѕ@������������������������       ���'�# @A            @Y@                           @�L���@�             s@������������������������       ���8@_            `b@������������������������       ����M�@g            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@      �@      ?@     �P@     `|@     �R@      �@      h@     ��@     0u@     �@@      �?     �T@     �e@      @      $@     �Z@      @     @}@     �E@     `q@      S@      @              8@     �L@                     �A@             `o@      *@     �`@     �@@                      1@      ;@                      <@             �R@       @      R@      :@                      &@      0@                      :@              J@      @      C@      6@                      @      &@                       @              7@      �?      A@      @                      @      >@                      @              f@      @      O@      @                      @      3@                                     �X@      �?      7@      @                      @      &@                      @             @S@      @     �C@       @              �?      M@     �\@      @      $@     �Q@      @      k@      >@      b@     �E@      @      �?      L@     �Z@      @      @     �M@      @     �i@      5@     �`@      >@      @      �?      @@     �F@      �?       @      @@      �?      J@      .@     @P@      0@      @              8@     �N@      @      @      ;@      @      c@      @     �Q@      ,@                       @      "@              @      (@              *@      "@      "@      *@      �?               @      @              @      (@              @      @      @      $@      �?                       @                                      "@       @      @      @              3@     �h@     @y@      ;@      L@     �u@     �Q@     ��@     �b@     Ѐ@     pp@      <@      3@      b@     �n@      4@      C@     �m@     �K@     �m@     �^@     `m@     `f@      9@      (@      G@     �Z@      "@      ,@     �U@      1@      M@     �D@      O@     �Q@       @       @      �?      2@      �?              3@      @       @      @      "@      6@              @     �F@     @V@       @      ,@      Q@      *@      L@      A@     �J@     �H@       @      @     �X@     @a@      &@      8@      c@      C@     `f@     @T@     �e@      [@      1@      @     �J@     �K@       @      1@     @R@      7@      \@      D@     @W@      N@      "@      @      G@     �T@      @      @     �S@      .@     �P@     �D@      T@      H@       @             �J@     �c@      @      2@     @[@      .@     pt@      ;@     �r@      U@      @             �C@     @[@      �?      @     �R@      @      q@      ,@     �j@      L@      @             �B@      Z@      �?      @     �L@      @     `n@      ,@     �e@     �K@       @               @      @                      2@      �?      ?@              E@      �?      �?              ,@      I@      @      &@      A@       @     �J@      *@     @V@      <@                      (@      @@      @      �?      $@      @      :@      @      E@      $@                       @      2@      @      $@      8@      @      ;@      @     �G@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ� F'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�i���$@�	           ��@       	                   �8@��'
\5@           `�@                           �?����6@{           ��@                            �?��Qؑ@R           ��@������������������������       ��(K�@S             a@������������������������       �ǿw @�            �x@                          �7@nx<�Fc@)           �}@������������������������       �9���"@           p{@������������������������       �/��U@             B@
                            @��8/H�@�             m@                          �<@Qϥ��@p             e@������������������������       ���F��@H            �Z@������������������������       ��Z*0�&@(             O@                           @��F�%@.             P@������������������������       ���Go-@'             J@������������������������       �|%��b�?             (@                           @���W�@�           �@                          �5@�p����@o           d�@                           @aV�,Uk@g           ��@������������������������       �"�M��@P           �@������������������������       ���-�@           P|@                           @v����@           @�@������������������������       ���KCO	@�           @�@������������������������       �5y�d+@           �z@                           �?;�}%g�@*            �O@������������������������       ��xb嫯@             2@                           6@�
�m0�@            �F@������������������������       �\<����@	             (@������������������������       ��5k��@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        (@     @r@     ��@      :@      K@     @|@     �U@     D�@      k@     0�@     @v@      ;@             �T@     `d@       @      &@      Z@      $@     �}@      D@     q@     �S@      @             �L@     @a@       @      "@     @T@      @     @z@      :@     �k@     �H@      @             �@@      S@       @       @     �I@      @     �l@      2@     @W@      2@      �?               @      2@              @      2@      �?     �P@              9@      @                      ?@      M@       @      @     �@@       @     �d@      2@      Q@      .@      �?              8@      O@              �?      >@             �g@       @     �_@      ?@       @              8@      K@              �?      >@             `f@      @      ]@      >@      �?                       @                                      &@      @      &@      �?      �?              9@      9@               @      7@      @      J@      ,@     �J@      >@      �?              .@      7@                      0@      @      ?@      @      E@      :@      �?              $@      *@                      $@      @      5@       @     �B@      @                      @      $@                      @      �?      $@      @      @      3@      �?              $@       @               @      @              5@      @      &@      @                      $@       @               @      @              *@      @      @      @                                                                       @              @                      (@     @j@     �y@      8@     �E@     �u@     @S@     ȁ@      f@     P@     Pq@      7@       @      i@     @y@      8@     �E@      u@     �R@     ��@     �d@      @     q@      5@      �?     �S@     @j@      @      :@     �b@      =@     Px@      O@     @s@     @[@      (@      �?     �H@     �`@      @      2@     �]@      5@     �m@      A@     `k@     �T@      @              =@     �S@      �?       @      ?@       @     �b@      <@     @V@      :@      @      @     �^@     @h@      4@      1@     @g@      G@     �e@      Z@     �g@     �d@      "@      @     @U@     �a@      ,@      *@      `@      C@     �S@     �T@     �X@      ]@      "@      �?      C@      K@      @      @     �L@       @     �W@      6@      W@      H@              @      "@       @                      (@       @       @      &@      @      @       @      @      �?      @                      @                       @              @       @               @      @                      "@       @       @      "@      @      �?                              @                       @      �?      @              �?      �?                       @       @                      @      �?      @      "@       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJj�)RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@h��K�g@�	           ��@       	                     @ ���d@F           �@                           �?��AYD@W           �@                           �?>8+�h�@�           ��@������������������������       �S�=�@�            �x@������������������������       ���p�o	@�            �v@                           @�]�A��@�           8�@������������������������       ��K��@�           h�@������������������������       ��wQ�W]@�           �@
                          �3@GΝ�;.@�           �@                           @��-X��@�            �v@������������������������       �ӽD��~@�            u@������������������������       �      @             8@                           @����:@           �y@������������������������       ����P�@�             t@������������������������       ��|@?            @V@                           �?���aI	@N           ؍@                           �?gGJ�f\@�            �p@                          @@@�"�P�Y@Z             c@������������������������       �E��@��@S            @a@������������������������       �%��,��?             ,@                          �:@��]�@@             \@������������������������       �"� ��,�?             F@������������������������       �x�f:�@%             Q@                           @,.?�	@�           ��@                           @�b0���	@,            ~@������������������������       �o�T�@A             Z@������������������������       �3�.�	@�            �w@                          �:@�'�j2D@�            `j@������������������������       ��+V�V@7            �S@������������������������       �R��@Q            �`@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B�        &@     pr@     `�@      B@     �P@     ~@     @S@     p�@      g@     ��@     @y@     �C@      @     �i@      z@      7@     �E@     Pv@     �B@     h�@     �Y@     �@     �o@      ;@      @     @c@     �s@      ,@      A@     p@      8@     (�@      S@     `|@     `d@      (@             �K@     @Z@       @       @     �P@      @     �s@      2@     @d@      ;@      @              ;@      J@       @       @     �C@      @     @d@      .@     @R@      (@       @              <@     �J@                      ;@             �b@      @     @V@      .@      �?      @     �X@     �j@      (@      :@     �g@      1@     �v@      M@     @r@      a@      "@      @      K@     �V@      $@      2@      ^@      "@     @Z@      H@      Z@     �T@       @       @     �F@     �^@       @       @     �Q@       @     0p@      $@     �g@     �J@      �?      �?      J@     @Y@      "@      "@      Y@      *@      i@      :@     `c@     @V@      .@              5@     �E@              @     �@@      @     �_@      &@     �P@      J@                      5@      D@              @      8@      @      _@      "@      O@     �H@                              @                      "@      �?       @       @      @      @              �?      ?@      M@      "@      @     �P@       @     �R@      .@     @V@     �B@      .@      �?      <@      I@      "@      @      M@      @      C@      .@      Q@      =@      (@              @       @                      "@      �?      B@              5@       @      @      @     @V@     @a@      *@      8@      _@      D@      `@     �T@     `b@      c@      (@              8@     �C@              @      ?@      @      K@      *@      I@      D@       @              7@      :@              @      6@      �?      1@      @      2@      @@       @              7@      7@               @      .@      �?      1@      @      1@      @@       @                      @              @      @                              �?                              �?      *@                      "@      @     �B@      @      @@       @                                                      �?      @      3@              ,@      @                      �?      *@                       @              2@      @      2@      @              @     @P@     �X@      *@      3@     @W@      A@     �R@     �Q@     @X@      \@      $@      @      B@     �R@      "@      0@      Q@     �@@      B@      L@     �I@     �U@      $@      @      $@      6@      �?      @      (@      @              1@      "@      0@      @              :@     �J@       @      *@      L@      <@      B@     �C@      E@     �Q@      @              =@      8@      @      @      9@      �?     �C@      ,@      G@      :@                      @      $@      �?      �?      @              2@      $@      2@      $@                      9@      ,@      @       @      2@      �?      5@      @      <@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJDz�IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?U�y�_j@�	           ��@       	                    �?ܸ���@           t�@                            �?R.��1�@�           ��@                           �?Ƣ��O@d             c@������������������������       �x1?�@'            �N@������������������������       ��A��/�?=             W@                            �?�3�;@C           �@������������������������       ��\���@|            �i@������������������������       ��Q�u�B@�            �r@
                           �?��N��@h           H�@                            @�/��a�@�            �n@������������������������       ��t�=1n@_            `b@������������������������       �f��,M�@;            �X@                           @VV��5�@�            0u@������������������������       ��?'$��@\            �b@������������������������       �G���b@r            �g@                           @Q�ws;@�           ؤ@                          �7@*w�f��@�           �@                           @ �M�@�           ��@������������������������       �D1L~��@�           ԑ@������������������������       �"{
 �@           �z@                          �;@Y�_I��	@�           h�@������������������������       ��[����@           �{@������������������������       ���5�	@�            Ps@                           @�z��	@�            �u@                           �?vM�Ω	@�            `i@������������������������       ��̇��	@^            �b@������������������������       ���SFd@%            �K@                          �4@��=��@\            `b@������������������������       �0��ƫ�@%            �O@������������������������       �ҍ&P*A@7             U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@      s@     �@      B@      L@     `|@     �V@     (�@     �i@     Ȉ@     �u@     �B@       @     @V@      f@      @      "@     �Y@      .@     �{@     �D@     �p@     @U@      @       @      C@     �W@      @      @      L@      &@     `p@      9@     @\@     �G@               @       @      ;@              �?      &@      @      Q@       @      ?@      @               @       @      0@                       @      @      *@       @      *@       @                              &@              �?      @             �K@              2@      @                      B@     �P@      @      @     �F@       @     @h@      7@     �T@     �D@                      3@      =@       @      �?      5@      @     �P@      $@      9@      <@                      1@      C@      @      @      8@      @     �_@      *@     �L@      *@                     �I@     �T@      �?       @     �G@      @     �f@      0@     `c@      C@      @              <@      G@               @      ?@              H@      "@     �G@      =@      @              0@      .@               @      5@              <@      @      C@      2@      @              (@      ?@                      $@              4@      @      "@      &@                      7@      B@      �?              0@      @     �`@      @      [@      "@      �?              ,@      1@                      &@      �?      K@      @     �H@              �?              "@      3@      �?              @      @      T@      @     �M@      "@              (@      k@     �x@      >@     �G@     �u@      S@     H�@     �d@     h�@     �p@      >@       @     �f@     �u@      9@     �E@     0s@      P@     0~@     �_@     `~@     �l@      1@       @      ]@     Pp@      $@      5@      h@      ?@     x@     �Q@      v@     @^@      @       @     �W@     �e@      @      *@     �b@      >@     �p@      D@     �p@     �W@      @              5@     @V@      @       @     �F@      �?     �]@      ?@      U@      :@      �?      @     �P@      V@      .@      6@     �\@     �@@     �X@     �K@     �`@     �Z@      &@      �?     �A@     �G@      $@      &@     �Q@      $@      P@      B@     �W@      J@      "@      @      ?@     �D@      @      &@     �E@      7@      A@      3@      D@     �K@       @      @     �A@      H@      @      @      F@      (@     �Q@      C@     �C@      C@      *@      @      6@      A@      @      @      ?@      $@      ;@     �@@      "@      4@      @      @      .@      4@      @       @      <@      @      5@      3@      @      1@      @              @      ,@              �?      @      @      @      ,@      @      @                      *@      ,@       @      �?      *@       @     �E@      @      >@      2@      @              @      @              �?      �?              8@              .@      *@                      $@       @       @              (@       @      3@      @      .@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�"EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?S���ZB@�	           ��@       	                    @h`�a@O           �@                           �?��1�{�@3           ��@                           �?-uQ�@�            @s@������������������������       ���z��@:            �U@������������������������       �EDs��@�            �k@                            �?Lf/>	@h            �@������������������������       �B�fЖ�@�            pr@������������������������       ��g��@�            �q@
                          �4@��4@           p�@                          �1@��އ@5           �}@������������������������       ���?N@v            �f@������������������������       �0zBp��@�            pr@                           @��0��r@�             w@������������������������       ��e�6�@�            �o@������������������������       ����Z0�@J            �\@                           @$:���N@h           �@                           �?p�ǔV�@d           P�@                           �?���O
	@�           p�@������������������������       ����x�@�            �w@������������������������       �>L�y)�	@�           ��@                          �2@
P>K�@�            `v@������������������������       �'�`���@:            @W@������������������������       �����g+@�            �p@                            @q[��j@           ��@                           @Q�����@�           Є@������������������������       �]fZ��9@           �|@������������������������       ���4�J�@�             j@                           @q��Q,@]             c@������������������������       ��b�2���?B            �Z@������������������������       ���E�a@             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     @s@     ؁@      1@     @Q@     �{@     �Q@     `�@     �m@     ؈@     �u@      <@      @      ^@      q@      "@      ;@      i@      C@     �}@     @\@     �s@      b@      "@      @      S@     @a@       @      4@     �^@      @@      e@     @W@     �]@     @X@      @              6@      D@      �?      $@      B@      @     �U@      7@      K@      >@      �?              @       @                      &@              <@      @      <@      @                      3@      @@      �?      $@      9@      @      M@      3@      :@      :@      �?      @      K@     �X@      @      $@     �U@      ;@     �T@     �Q@     @P@     �P@      @              2@      L@       @       @      E@      3@      @@      J@      >@      ?@      @      @      B@      E@      @       @      F@       @      I@      2@     �A@      B@               @      F@     �`@      �?      @     �S@      @      s@      4@     �h@      H@      @              4@     �Q@      �?      @      >@              i@      (@      \@      :@                      @      9@              @      (@              V@      �?     �D@      @                      ,@      G@      �?              2@             @\@      &@     �Q@      5@               @      8@     �O@               @     �H@      @     @Z@       @      U@      6@      @       @      0@     �D@                     �@@      @     @V@      @      I@      *@      @               @      6@               @      0@       @      0@      @      A@      "@              (@     �g@     �r@       @      E@     `n@     �@@     ��@      _@      ~@     �i@      3@      (@      b@     �h@       @     �@@     �g@      <@     @l@      Y@     `o@     �c@      1@      (@     @[@     �a@      @      ;@     @b@      7@     @a@     �R@     `g@     �_@      1@      �?      @@     �O@       @      @      F@      @     �P@      5@      S@      K@      @      &@     @S@     �S@      @      5@     �Y@      0@      R@     �J@     �[@      R@      *@              B@      M@       @      @     �E@      @      V@      :@      P@      >@                      @       @               @      @       @     �D@      @      1@      (@                     �@@      I@       @      @      D@      @     �G@      5@     �G@      2@                     �E@      Y@              "@      K@      @      s@      8@     �l@     �H@       @              ?@     @W@              @     �E@      @     �n@      6@     `f@     �E@       @              2@     @Q@              @      <@      �?     `g@      $@     �]@      7@                      *@      8@               @      .@      @     �L@      (@      N@      4@       @              (@      @              @      &@      �?      N@       @      I@      @                      @      @                      @      �?      G@       @      D@      @                       @      @              @      @              ,@              $@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJꇣDhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @f�0��G@�	           ��@       	                    �?��s+��@�           z�@                           �?ǬIS��@�           @�@                           �?�"[0�@�            `t@������������������������       ��M�$!@.            �Q@������������������������       �D��=@�            �o@                          �7@Ě-���@�             v@������������������������       ������@�            `n@������������������������       ��L'׶@B            �[@
                           @��%!Q	@�           T�@                           �?
��]$	@�           h�@������������������������       ���7M�	@�           T�@������������������������       �����b@�            Px@                          �8@3[1BW@#            �M@������������������������       �"��A��@            �D@������������������������       �D�9�<@
             2@                          �4@��z��@:           0�@                           �?���@O           ��@                          �0@��2O���?�            �v@������������������������       ������?#            @P@������������������������       ���"���?�            �r@                           @�3���T@l           �@������������������������       ��$�\�@W            @`@������������������������       �=��/)`@            z@                          �5@����l@�           ��@                           @X�z@f            `c@������������������������       �jŉҨ@_             b@������������������������       �QcX^@             $@                           @��a�@�           �@������������������������       �z���R@z           ��@������������������������       �xC��� @             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pr@     �@      D@     �J@     �|@     �Q@     ��@      k@     ��@      w@      ?@      1@     �j@     �s@      ?@     �C@     �t@     �I@     Px@     �f@     �w@      p@      ;@      @     �R@      Y@       @      "@     @Q@      @     @f@      C@     �a@      L@      @      @      D@     �D@       @      @     �A@      @      Y@      0@     �H@      =@      �?      @      @      "@                       @              <@              .@      @                     �A@      @@       @      @      ;@      @      R@      0@      A@      :@      �?             �A@     �M@               @      A@             �S@      6@     @W@      ;@      @              <@      @@              �?      6@             �N@      (@     �Q@      1@                      @      ;@              �?      (@              1@      $@      7@      $@      @      ,@      a@     `k@      =@      >@     Pp@      H@     `j@      b@      n@      i@      6@       @      `@     �j@      =@      >@      o@     �G@     @j@      a@      m@     �h@      1@       @      \@      c@      7@      7@     �f@     �C@     @`@     �Z@     �d@     `b@      1@              1@     �N@      @      @     �P@       @      T@      =@     @P@      I@              @       @      @                      (@      �?      �?      "@      "@      @      @      @       @      @                      "@              �?      @      @      @      @      @               @                      @      �?              @      @                      �?     @T@     @l@      "@      ,@     �_@      3@     Ѓ@      A@      z@      \@      @              G@     �\@      @      "@     �H@      @     �z@      .@     �i@     �E@                      &@     �B@               @      ,@             @i@      @      T@      ,@                              ,@                      @             �@@              @      @                      &@      7@               @       @              e@      @     �R@       @                     �A@     @S@      @      @     �A@      @     �k@      "@      _@      =@                      2@      ;@                      &@       @      E@      @      2@       @                      1@      I@      @      @      8@      �?     �f@      @     �Z@      5@              �?     �A@      \@      @      @     @S@      0@      j@      3@     �j@     @Q@      @              �?      B@                      "@      @     �D@              J@      @      @              �?      B@                      "@      @      D@             �H@      @       @                                                      �?      �?              @      @       @      �?      A@      S@      @      @      Q@      $@      e@      3@      d@     �O@              �?      >@      S@      @      @     �O@      "@     �d@      .@      d@     �O@                      @                              @      �?      �?      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJF�rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@���j�T@�	           ��@       	                    @��i��@�           ��@                           �?� ���@+            ~@                           �?�j~N@y            �i@������������������������       ����ߠ�@4            �W@������������������������       �`x^�@E            �[@                           �?�^t�4z@�            0q@������������������������       ���c�@             2@������������������������       �b:�T@�            p@
                           @��/?�� @Z           �@                           @/^*&��?�            �y@������������������������       ��`��|>�?=            �X@������������������������       �;��"M��?�            �s@                           @��'4�@f            �d@������������������������       �p�����?             L@������������������������       ��C2$�C@G            @[@                           @�6g�4@           N�@                           �?J)2f	@/           \�@                           @{�zН�	@           ��@������������������������       �r���n�	@�           ��@������������������������       �k$>U_	@M            �]@                           @ю<��@            {@������������������������       ��<e�G@�            �w@������������������������       ���滉�@!            �I@                            �?C(�B@�           @�@                           �?0�K>	@�            �@������������������������       ��f�� @s             g@������������������������       �����%@           �z@                          �7@/(տ�D@V           `�@������������������������       �Š�&�@�            �t@������������������������       �[D�T�@�            @l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �s@     (�@      5@     �F@     �}@      W@     8�@      m@     P�@      u@     �B@      �?     �H@      _@      �?      @      [@      @     0z@      L@     �k@      Q@       @      �?      9@      L@      �?       @      U@      @     @`@      G@      U@      H@                       @      9@                      =@      @     �Q@      ,@      F@      &@                      @      ,@                      4@      @      >@      $@      "@       @                      �?      &@                      "@             �D@      @     �A@      "@              �?      1@      ?@      �?       @     �K@             �M@      @@      D@     �B@                               @              �?      @              �?      @              @              �?      1@      =@      �?      �?      I@              M@      ;@      D@     �@@                      8@      Q@              @      8@             r@      $@      a@      4@       @              6@      H@                      1@             �l@      @     �T@      @       @              @      8@                      �?              O@              "@                              3@      8@                      0@              e@      @     @R@      @       @               @      4@              @      @             �M@      @     �K@      .@                              @              �?      @              *@              =@      @                       @      ,@              @      @              G@      @      :@      (@              6@     �p@     �x@      4@     �C@     �v@     @V@     X�@      f@     h�@     �p@     �A@      4@     �g@     �o@      1@      >@     �m@      P@      o@      a@     0p@     �h@      ?@      4@     `b@     �g@      1@      9@      f@      J@      c@     �Y@     �g@     @c@      <@      .@     @a@     @e@      0@      9@     `d@      F@     @a@     @S@      g@      b@      4@      @      "@      3@      �?              *@       @      .@      :@      @      "@       @             �E@     @P@              @     �O@      (@     �W@     �@@     �Q@     �F@      @             �A@      J@              @      N@      (@     �V@      4@      P@     �D@      @               @      *@                      @              @      *@      @      @               @      T@     `a@      @      "@     @_@      9@     0w@     �D@     �r@     �Q@      @             �C@      V@               @     �P@      0@     �f@      4@     `c@     �D@      �?              �?      ;@                      ,@      @      T@      @      J@      @                      C@     �N@               @     �J@      *@     �Y@      0@     �Y@     �B@      �?       @     �D@     �I@      @      @      M@      "@     �g@      5@     �a@      >@      @              <@     �C@      �?              =@      "@      ^@      @      T@      3@       @       @      *@      (@       @      @      =@              Q@      2@     �O@      &@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�3s|hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�4�.@�	           ��@       	                    �?�UM�xj@           �@                            @�'��@4            @                          �;@4o
{�"@�            �q@������������������������       ���M�^�@�            �n@������������������������       �j�F��@            �C@                          �<@N�c�1�@x            �j@������������������������       ���l��6@n            �h@������������������������       �>��_�@
             0@
                          �2@�.�P.@�           ��@                          �0@Ɵ�*d	�?�            �r@������������������������       ��k�^%�?*            �R@������������������������       �e�P�>�?�            �k@                           �?��@�H@,           �~@������������������������       �,^�fv�@�             q@������������������������       �H���@�            @k@                          �4@+_��
@�           ��@                           �?gm#~�A@�           ��@                          �3@&m��T4@>           �~@������������������������       �@u�Ą@�            `w@������������������������       ��/�Z��@I             ]@                           @���V@�           ȅ@������������������������       ��S`֝�@�           �@������������������������       �n�Bf�@             8@                            �?.�T�V	@�           ��@                           @Ь~,Z2	@�             y@������������������������       �~�rt>�	@�            pq@������������������������       �|�ք�@M            �^@                          �:@�N�t��@�           @�@������������������������       �֎c@�           `�@������������������������       �����^�	@�            @r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     pq@     �@      6@     �N@     @|@      Q@     ��@     �m@     8�@     �v@      9@      �?      V@     �f@      @      @      Z@      @     `z@     �F@     �t@     �U@      @      �?      K@      S@      @      @     �L@      �?     �[@      =@     �[@     �F@      @      �?      >@      G@              �?     �A@              I@      .@     �R@      ;@      @              :@      E@              �?      =@              H@      (@     �P@      0@      @      �?      @      @                      @               @      @       @      &@                      8@      >@      @      @      6@      �?      N@      ,@      B@      2@                      7@      :@      @       @      2@      �?      N@      (@     �A@      1@                      �?      @              @      @                       @      �?      �?                      A@     �Z@                     �G@      @     �s@      0@      l@      E@      �?              &@      A@                      &@             @c@      �?     �Q@      .@                              1@                      @              B@              *@      @                      &@      1@                      @             �]@      �?     �L@      (@                      7@     @R@                      B@      @     �c@      .@     @c@      ;@      �?              (@     �D@                      7@      @     @Y@      ,@      O@      1@                      &@      @@                      *@      �?     �L@      �?      W@      $@      �?      ,@     �g@     `v@      3@     �K@     �u@      O@     P�@     @h@     ��@     Pq@      5@      @     �J@      c@      @      (@     @c@      (@     �t@     �P@     �p@     �]@      "@      �?      .@      S@      @      @     �R@      @     @_@     �@@      Y@     �I@              �?      .@     �N@      �?      @     �J@       @     @Z@      6@     �S@     �@@                              .@      @      @      5@      @      4@      &@      6@      2@              @      C@      S@      @      @      T@      @      j@     �@@     �d@     �P@      "@      @      B@      S@      @      @     @R@      @     �i@     �@@     �c@     �P@      @               @                              @       @       @              @      �?      @      $@     @a@     �i@      (@     �E@     @h@      I@     �k@      `@     �p@     �c@      (@      @     �I@      F@      @      *@     �G@      $@      Q@      H@     �L@     �J@       @      @      C@      =@       @      *@     �C@       @      B@      E@      =@      B@       @              *@      .@       @               @       @      @@      @      <@      1@              @     �U@     @d@       @      >@     `b@      D@      c@      T@     �j@     �Z@      $@      @     �N@     �a@      @      2@     �Y@      6@     @\@     �G@     `d@      Q@      @       @      :@      6@      @      (@     �F@      2@     �C@     �@@      I@      C@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�M�0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���b�T@�	           ��@       	                    @yK�\A@�           ��@                           �?�"C�-X@?           ��@                          �3@�t\�@�            `u@������������������������       ���Y�y@�            pp@������������������������       ��g�ҡ@5            �S@                           �?�5�s�@b           �@������������������������       ��X<O�@m            �e@������������������������       �A1��A�@�            Pw@
                           �?�L����@H           h�@                            �?����>��?�            �v@������������������������       ��Ҝ��7�?:            @X@������������������������       ����ʓ @�            �p@                            �?ʹ�u�8@]           ��@������������������������       �#�)W�@�            �v@������������������������       �Z�8~@�             j@                           �?�(���@            H�@                           �?]H�&�V@}            �@                            �?��`�t@�            �r@������������������������       ���q�)1@n            �f@������������������������       ��r-���@O            �\@                            �?.Ը^�@�            �s@������������������������       ���7���@*             R@������������������������       ��1�FrJ@�            @n@                            �?Q�	�0	@�            �@                          �<@"�ŕ	@�           Ȉ@������������������������       �.1�L�	@�            �@������������������������       �RW�A�@N            @^@                           @�V�K�z@�           8�@������������������������       ��"�R1@`            �c@������������������������       ��Y�X@Q           X�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     ps@     �@     �A@     �L@      @     �S@      �@     �j@     ��@     �w@      6@       @     �[@     @j@      &@      1@      g@      ,@     ��@     �V@      y@      c@      @       @     �O@     @[@      "@      @      a@      (@     �i@      S@      e@      X@      @              1@     �L@      @      �?     �J@      @      U@      B@      E@     �C@       @              "@      H@      �?             �B@      @     @Q@      8@     �B@     �@@      �?               @      "@      @      �?      0@              .@      (@      @      @      �?       @      G@      J@       @      @     �T@       @     @^@      D@     �_@     �L@      @              3@      4@                      3@              J@      @     �H@      &@               @      ;@      @@       @      @      P@       @     @Q@     �B@     @S@      G@      @             �G@     @Y@       @      $@     �H@       @     �z@      ,@      m@      L@      �?              &@      @@              @      *@             �j@      @     @R@      *@      �?                      $@                      �?             �Q@              (@      @                      &@      6@              @      (@             �a@      @     �N@      $@      �?              B@     @Q@       @      @      B@       @     �j@      "@     �c@     �E@                      .@      D@       @      @      ;@             �`@      @      \@      ?@                      5@      =@               @      "@       @     @T@      @     �G@      (@              2@      i@     �r@      8@      D@     ps@      P@      y@     @_@     �v@     �l@      0@       @      N@     �W@      @       @     @R@      @     @d@      5@      a@     �E@       @       @     �C@      G@      �?       @      H@      �?     �G@      .@      N@      >@      �?       @      8@      7@              @      ;@      �?      :@       @     �E@      9@      �?              .@      7@      �?      @      5@              5@      @      1@      @                      5@      H@      @              9@      @     �\@      @      S@      *@      �?                      *@      @              @      @     �@@               @      @      �?              5@     �A@                      2@       @     �T@      @      Q@      $@              0@     �a@     @i@      4@      @@     �m@     �L@     �m@      Z@      l@     @g@      ,@      *@     �S@     @Z@       @      3@     @\@     �C@     �]@     �Q@     @\@     �Z@      @      (@      P@     �V@       @      3@     @X@      =@     �\@     �J@     �Z@      R@      @      �?      .@      ,@                      0@      $@      @      2@      @     �A@      �?      @      O@     @X@      (@      *@     @_@      2@     �]@     �@@     �[@     �S@      @       @      &@      ;@       @       @      C@      @      @      (@     �A@      .@              �?     �I@     �Q@      $@      &@     �U@      *@      \@      5@      S@      P@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ7��chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @ w�\@�	           ��@       	                     �?1�b�@�           ��@                          �4@L��J��@�           ��@                          �2@?���C�@�            �q@������������������������       �}a>"#�@[            @c@������������������������       ��QuOLh@G            �`@                          �:@����
@           @{@������������������������       ��K 
@�            �s@������������������������       �@�9��@J            �]@
                            @P|�a�@�           �@                          �4@�r�'	@�           ��@������������������������       �ب#�L�@�            @s@������������������������       � ����	@           �x@                           @l��]�@           0�@������������������������       �Hd��=@�           ��@������������������������       ��,b���@�            �i@                           �?�x��k�@)           ԙ@                            @�y m.� @a           X�@                          �4@⫒�x@&           �|@������������������������       ��!�:��?�            �r@������������������������       �p8���@o            �d@                           7@��P��?;            �W@������������������������       ����,�j�?3            @T@������������������������       ��!�S�0�?             ,@                            �?�XV�@�           (�@                           �?�r8���@�            �n@������������������������       ����z�@L            @[@������������������������       ��C�Z @U            �`@                           @�D�qq{@'           ��@������������������������       ��%��k6@�           Ȃ@������������������������       �̆k_X@�            �o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     �@      <@     @P@     p}@      Y@     H�@     �k@     �@      u@     �@@      0@     `j@     �s@      4@      K@     Pu@     @T@      z@     @e@      w@     �m@      <@      @     �K@     �U@      @      1@      [@      9@     �c@      O@      _@      O@      0@              .@      8@                     �F@       @     �X@      7@      L@      3@      @              @      3@                      0@       @     �O@      @     �A@      @                      "@      @                      =@              B@      1@      5@      (@      @      @      D@      O@      @      1@     �O@      7@      N@     �C@      Q@     �E@      *@      @      A@      I@      @      1@      B@      *@      J@      >@      G@      8@      $@              @      (@       @              ;@      $@       @      "@      6@      3@      @      *@     �c@     �l@      .@     �B@      m@      L@     p@      [@     �n@      f@      (@      @      U@     @T@      @      0@     @Z@      9@     @]@     �I@     �[@     @V@       @       @      =@      =@      @       @      K@      @     �R@      3@     �P@      ;@              @     �K@      J@      @      ,@     �I@      6@     �E@      @@     �F@      O@       @      @      R@     �b@       @      5@      `@      ?@     �a@     �L@     �`@     �U@      @      @      K@      Z@       @      *@     �Z@      0@     @]@     �@@      [@     �O@      @      @      2@      G@               @      5@      .@      7@      8@      9@      8@              �?      S@     @h@       @      &@     @`@      3@     ��@      J@     {@     �X@      @              $@     �P@      �?      @     �B@      @     q@      $@     �`@      2@                      "@      P@      �?       @     �@@      @     `k@      @     �Z@      1@                       @      @@               @      (@              d@      @     @Q@      "@                      �?      @@      �?              5@      @      M@       @     �B@       @                      �?      @              �?      @              K@      @      :@      �?                              @              �?      @             �G@              9@      �?                      �?                                              @      @      �?                      �?     �P@     �_@      @       @     @W@      .@     v@      E@     �r@      T@      @              4@      1@      �?              .@             @Y@      &@     @P@      ,@                      @      (@                      &@              =@      @     �B@      $@                      ,@      @      �?              @              R@      @      <@      @              �?      G@     �[@      @       @     �S@      .@     �o@      ?@     �m@     �P@      @      �?      A@      Q@       @       @      I@       @      j@      6@      e@     �A@       @              (@      E@      @      @      <@      @     �E@      "@      Q@      ?@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJS�]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����@�	           ��@       	                     @uд���@�           L�@                           �?��H_�@l           T�@                           �?ŉd�
 @             }@������������������������       ��08T#@�            �k@������������������������       ��e��?�@�            �n@                            �?�	GdL@	@L           �@������������������������       ��Ș�us	@�           ��@������������������������       ��� �H@V            �a@
                          �1@�U3T@           ��@                          �0@�#X���@A            �W@������������������������       ��;�\�Z@             3@������������������������       ���*���@4             S@                          �9@��O�@�           ��@������������������������       ��L�C}�@\           ��@������������������������       ���eN��	@~            �g@                           @�Z{h�@1           ��@                            �?�L*�@�            0x@                           @�a�mԟ@@            �X@������������������������       ���U��@/            �Q@������������������������       ���F��@             ;@                           �?�,�q�@�            r@������������������������       �����t�@A            �Y@������������������������       ��0VtC�@x            @g@                           @����z�@8           ��@                            �?�F^�B@�            �@������������������������       ��4��M�@             y@������������������������       �Z�-?�% @�             w@                           �?aRŲ��@T           ��@������������������������       ��J��G�@�            0q@������������������������       �0zm=��@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     x�@      @@     �J@     p|@     �O@     \�@     @e@     ��@      v@      @@      2@     �k@     0u@      7@      F@      t@      F@     Px@     `a@      y@     �n@      ;@       @     �_@      h@      "@      :@     �h@     �B@     �m@      X@      o@      e@      1@      �?      E@     �K@      �?      @      J@      @      ]@      .@     �]@      K@      @      �?      2@      <@      �?      @      ;@      @      J@      (@      F@      >@                      8@      ;@                      9@      �?      P@      @     �R@      8@      @      @      U@     @a@       @      6@     `b@     �@@     �^@     @T@     @`@     �\@      *@      @      Q@      ^@       @      3@     @_@      ?@     @Y@      R@     �[@     �T@      *@              0@      2@              @      6@       @      5@      "@      3@      @@              $@     @X@     @b@      ,@      2@     �^@      @     �b@     �E@     @c@      S@      $@              @      &@       @              "@             �@@       @      6@      @                              @                      @              @      @      @                              @       @       @              @              >@      @      1@      @              $@     @W@     �`@      (@      2@     �\@      @     �]@     �A@     �`@     �Q@      $@      @      N@      \@       @      $@     �V@      @      W@      3@     �Z@     �H@      @      @     �@@      7@      @       @      8@      �?      :@      0@      :@      5@      @      �?     @S@     �k@      "@      "@     �`@      3@     ��@      ?@     �z@      [@      @      �?      :@      P@                      ?@      (@     �`@      $@      U@      8@      @              $@      $@                      @              C@      @      3@      &@                       @       @                      @             �A@      �?      *@      @                       @       @                                      @      @      @      @              �?      0@      K@                      :@      (@     �W@      @     @P@      *@      @               @      *@                      @       @     �G@       @      8@      �?              �?       @     �D@                      4@      $@     �G@      @     �D@      (@      @             �I@     �c@      "@      "@     �Y@      @     p�@      5@     �u@      U@       @              ;@     �V@      �?       @      I@       @     Pv@      "@      h@     �D@                      .@      M@      �?              :@       @     `e@       @     @Y@      4@                      (@      @@               @      8@             @g@      �?      W@      5@                      8@     �P@       @      @      J@      @      e@      (@      c@     �E@       @              .@      @@      @      @      7@      �?     @Y@      @     �O@      8@                      "@      A@      @      @      =@      @      Q@      @     @V@      3@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��:��@�	           ��@       	                    �?���u�@�           ��@                            �?�J�V}@�           0�@                          �;@��e�'@�            �l@������������������������       ������[@�             k@������������������������       �XL��J@
             *@                            @��:�� @$           ~@������������������������       �c� ��@�            @n@������������������������       ��r�f�@�            �m@
                           �?�"�9iX	@�           �@                           @S�E|�	@�           ��@������������������������       �M�{f�`	@z           ؎@������������������������       ���τ�@W             b@                           �?϶ĝ ~@           �y@������������������������       �`{5�[@             F@������������������������       ��֟���@�            �v@                          �7@;��4j0@%           ��@                           �?�����@           L�@                           @��O9�?           �z@������������������������       �Ⱦ�����?�            �r@������������������������       ����P޽ @T             `@                           @$��7@           8�@������������������������       ��ŉE:C@r            �f@������������������������       �K�{��@�           ��@                          �<@2zRl@�@           �z@                          �9@�uf�G@�             u@������������������������       �ɰ�1�@{            �g@������������������������       ����L�@_            `b@                            �?�d��v*@7             V@������������������������       ���	;�@             F@������������������������       ��3f��@             F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     0t@     ؁@      7@     �J@     0{@      Q@     ��@     @j@     �@     0u@      =@      :@     @m@     �u@      0@      D@      t@     �L@     x@     @f@     �w@      n@      ;@      �?     �N@     �S@      @      "@     �W@      @     @j@      @@     `c@     �K@      @      �?      0@     �@@              �?      <@      �?     �N@      @     @P@      *@      @              ,@      =@              �?      ;@      �?     �N@      @     @P@      $@      @      �?       @      @                      �?                                      @       @             �F@      G@      @       @     �P@       @     �b@      ;@     �V@      E@       @              ?@      5@      �?      @      C@       @      N@      0@      H@      4@       @              ,@      9@       @      @      =@             @V@      &@      E@      6@              9@     �e@     �p@      *@      ?@      l@      K@     �e@     @b@      l@      g@      4@      9@     `a@     �h@      *@      :@      f@      B@     �X@     @Z@     �b@      b@      4@      1@      `@     �d@      *@      :@     �b@      :@      V@     �U@     �a@     �`@      &@       @      $@      A@                      <@      $@      &@      2@      @      &@      "@              A@     @R@              @      H@      2@      S@     �D@      S@      D@                       @      @              @       @       @      @      @      @      @                      :@     �Q@                      D@      0@     @R@      B@     �Q@      B@                     @V@     �k@      @      *@     �\@      &@     H�@      @@     px@     �X@       @             �L@     �d@      @      @     �O@      @     ��@      2@     �q@     �L@       @              ,@     �F@       @              1@      �?      o@      @     �U@      @      �?              &@      <@                      $@      �?     `g@      @     �J@      @                      @      1@       @              @             �N@       @     �@@       @      �?             �E@     �^@      @      @      G@      @      t@      &@     �h@      I@      �?              (@     �@@                      @      @     �Q@      @      D@      &@                      ?@     @V@      @      @      D@      �?     @o@      @     �c@     �C@      �?              @@      K@       @      @      J@      @     @\@      ,@     �Z@      E@                      6@     �C@              @     �E@      @     �V@      ,@     @W@      =@                      .@      =@                      8@             �I@      @     �E@      6@                      @      $@              @      3@      @     �C@      @      I@      @                      $@      .@       @       @      "@      �?      7@              *@      *@                      @      *@                      @      �?      $@              �?       @                      @       @       @       @      @              *@              (@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?W���B@�	           ��@       	                    @vל��T@           ��@                          �<@����5@�           @�@                           �?&�}�~@           ��@������������������������       ��b�!@           p{@������������������������       ��&���@r             e@                            �?���IXK@-            @R@������������������������       �����G@             ,@������������������������       ����ӄL@%            �M@
                           @Ǣ8줹 @[           ��@                          �2@O!�ʖ/�?�            pw@������������������������       ��悖}�?^            @d@������������������������       ���)�.l@�            �j@                          �5@�l~b@v             i@������������������������       ����^I @K            �_@������������������������       �p�/2��@+            �R@                           @�D-�;@�           Ĥ@                           �?hI��fz	@�           x�@                          �9@�
v���	@�           �@������������������������       �*���3	@           @�@������������������������       ��yLJ#r
@�            �s@                           @��Y��@           �y@������������������������       �w�ǉ�@y            @h@������������������������       ���/4g�@�            @k@                           �?~}���@�           �@                          �6@�J� ��@.            @T@������������������������       ��t��|�@!             L@������������������������       ���;O@             9@                           @�sdѹ@�           ��@������������������������       �<ԛ@�           �@������������������������       �����P^@�            `q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      r@     ��@      8@     �L@     �|@     �V@     X�@     `i@     ��@     Pu@      =@             @T@     �e@       @      (@     @]@      ,@     @|@      ?@     pr@     �R@      @             �Q@      Y@      �?      "@     �T@      @     @e@      <@     �c@      J@      @             �O@     @U@      �?      @      R@      @     �d@      7@     �b@      ?@      @              G@     �Q@      �?      @      L@      @     @Z@      6@      Z@      8@      @              1@      .@              �?      0@       @      O@      �?     �G@      @                      @      .@              @      &@              @      @      @      5@      �?              @      @                      �?                               @      �?      �?              @      $@              @      $@              @      @      @      4@                      &@      R@      �?      @      A@       @     �q@      @     @a@      7@                      @     �B@                      :@      @     `i@      �?     �T@      *@                      @      $@                      @             �Z@             �@@      @                      @      ;@                      4@      @     @X@      �?     �H@      $@                      @     �A@      �?      @       @       @     �S@       @      L@      $@                      @      1@              @       @              P@      �?      >@      @                              2@      �?              @       @      .@      �?      :@      @              8@     �i@      y@      6@     �F@     �u@      S@     8�@     �e@     h�@     �p@      9@      7@     �b@     �o@      0@      ?@     `k@     �P@      k@      b@     �m@     �g@      6@      7@     �\@      f@      .@      6@     �e@     �K@     �`@     �X@     @f@     �a@      5@      &@     �V@     �_@       @      3@      b@      @@      Z@      M@     �a@      W@      &@      (@      8@     �H@      @      @      <@      7@      ?@     �D@     �A@     �I@      $@             �@@     @S@      �?      "@     �G@      &@     @T@      G@      N@      G@      �?              "@      :@              @     �@@      @      F@      ,@      C@      4@                      8@     �I@      �?      @      ,@      @     �B@      @@      6@      :@      �?      �?     �M@     `b@      @      ,@     �_@      $@     �t@      ;@     �q@     @S@      @      �?      @      0@               @      &@       @      &@      @      9@      �?                      �?      0@                      $@       @      @              3@      �?              �?      @                       @      �?              @      @      @                              J@     ``@      @      (@     �\@       @     @t@      6@     `p@      S@      @              :@      Y@               @     �T@       @     �p@      *@     �g@     �G@      @              :@      ?@      @      $@     �@@      @     �L@      "@     �Q@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?<�Ƌ�@�	           ��@       	                   �;@���e�p	@�           ��@                            @͊�r�	@Y           ��@                           �?�iC�R�@�           ��@������������������������       �}��uj@�            �v@������������������������       �j>g�,�	@           �z@                           �?��V��	@c           x�@������������������������       ��w�,J�@c            `e@������������������������       ���5���	@            @z@
                           �?��u�z	@�             o@                            @�;�z�/	@=            �W@������������������������       ��禭p�@#             N@������������������������       �P��}J@            �A@                          �<@:����@g            @c@������������������������       ��m����@             9@������������������������       �Pw�o@U             `@                          �4@K�^� 0@�           ҡ@                           �?��瑞M@�           4�@                            �?�!���@t           p�@������������������������       �,`7 �K@Z             a@������������������������       �[O�/Ͻ@           P|@                          �1@�?g��@�           ��@������������������������       ���:%�1 @�            �n@������������������������       �KΣ	�@�            �x@                           �?}Vv�ع@�           p�@                          �8@Iz��@�            �q@������������������������       ��ж־.@u             g@������������������������       ��}`t��@@            @Y@                           @�����_@�           ��@������������������������       ���1*7�@�           �@������������������������       ��n\��@L             _@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pr@     X�@      B@      N@      |@     �X@     ��@     �i@     ��@     px@      ?@      1@     @d@     @n@      2@     �D@      o@     �P@     �k@      `@     �o@     @j@      7@      @     �a@      j@      1@     �@@     �k@     �D@     �i@     �[@     �k@     @c@      5@      @      W@     �^@      "@      7@     �[@      0@     �_@      Q@     �\@     �X@      @              =@     �O@       @       @     �J@      @     �R@      9@      M@      G@      �?      @     �O@      N@      @      .@      M@      (@     �J@     �E@      L@     �J@      @      @      I@     �U@       @      $@     �[@      9@      T@     �E@     �Z@     �K@      ,@              *@      B@               @      6@      �?     �C@       @      A@      0@              @     �B@      I@       @       @      V@      8@     �D@     �A@      R@     �C@      ,@      $@      4@     �@@      �?       @      <@      :@      ,@      2@     �@@      L@       @      @      @      4@      �?      @      "@      (@      @      @      &@      1@              @      @      ,@      �?              @      @      @      @      @      ,@              @       @      @              @      @      @      �?              @      @              @      ,@      *@              @      3@      ,@      $@      *@      6@     �C@       @      @       @       @                      @      �?      @               @       @                      (@      &@              @      0@      *@      @      *@      4@      ?@       @      �?     ``@     �s@      2@      3@     �h@      @@     �@      S@     ��@     �f@       @             �H@     �d@      $@      &@     @R@      @     �~@      ?@     0s@     �U@      @              ;@     @Q@      @       @      H@             `l@      2@     �a@     �G@                      @      3@              �?      3@              H@       @     �@@      "@                      5@      I@      @      @      =@             `f@      0@      [@      C@                      6@      X@      @      @      9@      @     pp@      *@     �d@     �C@      @              @      :@                      @             �\@      @     @R@      .@      @              2@     �Q@      @      @      4@      @     �b@       @     @W@      8@              �?     �T@     �b@       @       @     �_@      <@      o@     �F@      p@     �W@      @              $@     �G@      @              1@      @     @Y@      @     @S@      1@      �?              @      :@      @              0@      @      S@             �G@      @                      @      5@                      �?       @      9@      @      >@      *@      �?      �?      R@     @Y@      @       @     @[@      5@     `b@      D@     �f@     �S@      @      �?      J@     @R@      �?       @      V@      .@      `@      >@      e@     �R@      @              4@      <@      @              5@      @      2@      $@      (@      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ"�bhhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�8)�*@�	           ��@       	                    @��N�aD@�           t�@                          �1@��:r��@1           ��@                           @)�
P�@�            @p@������������������������       � Dp@N            �`@������������������������       ��M�1�@Y            �_@                          �2@����I@�           ��@������������������������       ���u�@�            @l@������������������������       �7���@�             y@
                           �?�.��H�@[           (�@                           @$�`�v�?�            0v@������������������������       �{�U X��?;            �W@������������������������       ���o�U��?�            @p@                            �?Mg�l�O@t           �@������������������������       �g*g�/@�            0v@������������������������       �Qn�w@�            �k@                           @jg�A@,           X�@                           �?��aew.	@&            �@                           �?���=�@�             v@������������������������       �P?T>�?@�            @p@������������������������       ��� ��?@:             W@                          �<@�1ۚ�	@D            �@������������������������       ���8Q�$	@�           @�@������������������������       ��Nb7�	@q             g@                          �8@����O=@           `�@                           �?��*�:]@?           �@������������������������       ��:�z|^@�            Pp@������������������������       ����۩@�            �n@                           �?d�'���@�            s@������������������������       �HM�8L��?+            �L@������������������������       �*�S�=@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     �p@     @�@      9@     �N@     �|@     �U@     ��@     �k@     ��@     0x@      @@      @     �T@     �i@      $@      :@      f@      4@     ؄@      V@     �v@      e@       @      @      J@     �Y@      "@      (@     @\@      1@     �m@     �R@     �a@     @]@      @              $@      B@      �?       @      2@      �?     �W@      6@     �H@      :@                      @      *@                      *@              K@      0@      5@      ,@                      @      7@      �?       @      @      �?     �D@      @      <@      (@              @      E@     �P@       @      $@     �W@      0@     �a@     �J@     @W@     �V@      @              ,@      9@              @     �G@       @      K@      8@      ;@      <@              @      <@      E@       @      @      H@      ,@     @V@      =@     �P@     �O@      @              ?@     �Y@      �?      ,@     �O@      @     �z@      *@      l@     �I@      �?              (@      @@              @      1@              j@      �?     @R@      @      �?               @      *@                       @              F@              9@      @                      @      3@              @      .@             �d@      �?      H@      @      �?              3@     �Q@      �?      $@      G@      @     �k@      (@      c@      F@                      @      @@              @      <@             �a@       @     @Z@      :@                      (@      C@      �?      @      2@      @     �S@      @     �G@      2@              @     �g@     �s@      .@     �A@     �q@     �P@     Px@     �`@     0z@     `k@      8@      @     �a@     �i@      &@      :@     �f@      K@     @c@      _@     �i@      c@      1@      �?      @@      N@              @     �F@      @     @S@      .@     �S@      >@      @      �?      :@      J@              @     �C@      �?      B@      ,@     �L@      8@      @              @       @                      @       @     �D@      �?      6@      @              @     �[@     @b@      &@      4@     �`@     �I@     @S@     @[@      `@     �^@      *@      @     �V@     �`@       @      ,@     �]@      B@     �P@     �S@     �Z@     �T@      $@      @      4@      ,@      @      @      1@      .@      $@      ?@      6@      D@      @              G@     @[@      @      "@     @Y@      (@     `m@      $@     �j@     �P@      @              =@     �R@       @       @      K@      "@     �e@       @     @^@      @@      @              4@      I@               @      <@      @     �R@      �?      L@      1@      @              "@      9@       @              :@      @     �X@      �?     @P@      .@      �?              1@      A@       @      @     �G@      @     �N@       @     �V@     �A@                              @                              �?      7@      �?      6@      @                      1@      ;@       @      @     �G@       @      C@      @     @Q@      @@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�4���\@�	           ��@       	                    �?^ݱb@]           �@                           @�i����@�           ؅@                           �?�=zyD>@�            @x@������������������������       ���i��@r            �h@������������������������       �iߑ8�@}             h@                           �?�_)C�@�            ps@������������������������       �ph���j�?t             f@������������������������       ��Ț��*@R            �`@
                          �4@�8$[�N@�           �@                          �1@�V`��@�           ��@������������������������       ��:�y�7@�            @k@������������������������       ��2-���@           �y@                           @[�!\�V	@            �@������������������������       ��h��.�	@T           X�@������������������������       ��<�ް@�            �s@                           @���":@P           H�@                           �?���2�@�           P�@                           �?��f�@�           ��@������������������������       ������@�             k@������������������������       ������[	@^            �@                            @����k@�            �q@������������������������       �������@@            �\@������������������������       ���D�@p            @e@                            @��`��@�           ��@                           �?Y�5���@           �|@������������������������       ���e��@�            @k@������������������������       �ItM���@�            �m@                           �?�@M��I@�            �n@������������������������       �˃s?�?5            @S@������������������������       � ����@j             e@�t�b��
     h�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@      �@      ;@      N@     �|@     @W@     �@      k@     ��@      x@      7@      @     @e@     �q@      2@      B@     `j@     �M@     �@      _@     P{@     `l@      .@             �F@     @U@      @      @      J@      @     �o@      :@     `d@      L@      @             �B@     �J@      @      @      :@       @     �W@      7@     �Y@      C@      @              5@      5@      @      @      2@       @     �K@      5@      :@      7@      @              0@      @@                       @              D@       @     @S@      .@       @               @      @@       @              :@      @     �c@      @      N@      2@                      @      0@                      1@       @     @Y@              :@      "@                       @      0@       @              "@      �?      M@      @      A@      "@              @     @_@     @i@      *@     �@@     �c@      K@     0t@     �X@      q@     `e@      $@             �B@     @T@      @      @      N@      @     @h@     �A@     �`@     @R@      @              @      <@              �?      ,@      �?      U@       @     �I@      9@                      ?@     �J@      @      @      G@      @     �[@      ;@     �T@      H@      @      @      V@     @^@      @      =@     �X@      I@      `@     �O@     �a@     �X@      @      @     �K@     @Q@      @      8@     @S@     �D@     �L@      L@      Q@      O@      @             �@@      J@       @      @      6@      "@      R@      @     @R@      B@       @      (@     �`@     p@      "@      8@     �o@      A@     �{@      W@      t@     �c@       @      $@     @W@     �b@      @      5@      f@      =@     `g@     �S@      d@     �_@      @      $@     �R@     �[@      @      1@      a@      ;@      ]@      H@      [@      Y@      @              4@      >@              @      A@      @     �J@      &@      C@      5@              $@      K@     @T@      @      ,@     �Y@      5@     �O@     �B@     �Q@     �S@      @              3@      D@              @     �C@       @     �Q@      ?@      J@      :@                       @       @                      5@      �?      5@      .@      =@      &@                      &@      @@              @      2@      �?      I@      0@      7@      .@               @      D@     �Z@      @      @      S@      @     p@      *@     @d@     �@@       @       @      =@     �U@       @       @      K@      @      b@      "@     �W@      8@       @       @      ,@     �G@      �?       @      7@      �?     �Q@      @     �E@      $@      �?              .@      D@      �?              ?@      @     �R@      @      J@      ,@      �?              &@      3@      �?      �?      6@              \@      @     �P@      "@                      �?       @                      �?              J@      �?      2@       @                      $@      1@      �?      �?      5@              N@      @     �H@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJtŻ-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�CS� /@�	           ��@       	                   �;@�/����@           f�@                          �1@�+�_@�           �@                           �?�x����@�            `p@������������������������       �hτ�6�@G            �Y@������������������������       �%�#=��@c            �c@                          �3@i�aڮ@           ��@������������������������       �d�o.�@           Pz@������������������������       �w�!m��@           `�@
                            @�}���	@�             s@                           @��l�?	@t            �g@������������������������       �(���Õ@E            �]@������������������������       �FZ�Rb@/             R@                          �@@%�i��@I            �\@������������������������       ����
�K@B            @X@������������������������       ��>��l�?             1@                           �?��\D�@.           X�@                          �4@B��g� @n           �@                           @y݌��"�?�            w@������������������������       ��YV��?�            �p@������������������������       �u�Z���@H            �Y@                          �6@X؋+�@�             j@������������������������       ��?U��_@7            �T@������������������������       ���o$��@Q            �_@                           @�r8���@�           T�@                          �9@����-@{            �h@������������������������       ���Y��@j            �d@������������������������       �}N|��@             ?@                           @%t�nK�@E           ��@������������������������       ���Ҥ�@�           ��@������������������������       ����w�0@�            `n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      s@     ��@      7@      L@     �z@     @S@     0�@     �j@     ��@      x@      9@      7@      l@     �t@      0@     �H@     0r@      M@      y@     �e@     @w@     �p@      4@      &@     �g@     r@      ,@      D@     p@      F@     �w@      b@     @u@     @i@      1@       @      &@     �I@      �?      �?      ;@       @      V@      *@     �G@      3@               @      �?      8@      �?              ,@       @      >@      @      (@      &@                      $@      ;@              �?      *@              M@      @     �A@       @              "@      f@     �m@      *@     �C@     �l@      E@     r@     ``@     Pr@     �f@      1@      @      ?@      B@       @      @     �N@      $@     @W@     �@@      U@      M@      @      @     @b@     @i@      &@      @@      e@      @@     �h@     �X@      j@     @_@      ,@      (@     �B@     �E@       @      "@      A@      ,@      7@      <@      @@     �P@      @       @      2@      8@       @       @      5@      $@      (@      4@      ;@      F@       @      @       @      2@               @      &@      @      "@      @      .@     �@@       @      �?      $@      @       @              $@      @      @      ,@      (@      &@              @      3@      3@              @      *@      @      &@       @      @      7@      �?              0@      (@              @      $@      @      &@       @      @      7@      �?      @      @      @                      @                                                             �S@      j@      @      @     �a@      3@     ��@     �D@     �z@     @]@      @              *@     �P@              @     �A@      @     �r@       @      `@      8@                      &@     �C@              @      ,@             �j@      @     �Q@      *@                       @      ;@                      @             �d@      �?      J@      $@                      @      (@              @      $@             �H@      @      3@      @                       @      ;@                      5@      @     �T@      @     �L@      &@                              (@                      $@      @     �C@      �?      *@      @                       @      .@                      &@             �E@      @      F@       @                     �P@     �a@      @      @     @Z@      .@     @u@     �@@     �r@     @W@      @              (@      =@              @      1@      @     �L@      *@      D@      5@                      &@      :@               @      (@      @      L@      @      B@      (@                      �?      @              �?      @              �?      @      @      "@                      K@     @\@      @      �?      V@      &@     �q@      4@     0p@      R@      @             �B@     @U@                      O@       @     �l@      ,@     �g@     �D@      @              1@      <@      @      �?      :@      @     �K@      @      Q@      ?@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�S�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�앝�=@�	           ��@       	                    �?whP%�q@!           ��@                          �;@Z�,X�@1           �|@                          �2@�3���@            y@������������������������       ���G�o@G             Y@������������������������       ��nDPn@�            �r@                          �=@0A�/�=@$             L@������������������������       �:=I���@             9@������������������������       ��By��@             ?@
                            �?�_9':@�            �@                           @���+��@}             i@������������������������       �����n@>            �W@������������������������       ��_
���??            �Z@                          �7@Թp���@s           ؂@������������������������       ���~xT@#            }@������������������������       �hs�s�@P             a@                          �5@�ks5.@�           ��@                          �3@����ߛ@�           ,�@                           @�z�[��@;           ؋@������������������������       ��L�7@           p{@������������������������       �;�h@"           @|@                           @�m�b*:@K           ��@������������������������       �j���'@�            `o@������������������������       �4��b�@�            Pq@                           @(e�3H	@           H�@                           @�
���	@�           �@������������������������       �������	@�           ��@������������������������       ��,e�m�@?             \@                          �7@G�����@            {@������������������������       ��݈|o@[             b@������������������������       �d�[)\Q@�             r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     p�@      <@      M@     �|@      T@     @�@     �m@     ��@     �t@     �@@             @S@     @c@       @      @     �[@      *@     �}@     �G@     �p@      X@       @              F@     �Q@              @     �N@      �?     �X@      @@      W@      H@      @             �B@      N@              @      K@             @X@      <@     �U@      ?@      @              �?      (@              �?      $@              C@      @      5@      &@                      B@      H@               @      F@             �M@      6@     @P@      4@      @              @      $@               @      @      �?       @      @      @      1@                      @      @                      @      �?               @       @      @                      @      @               @      @               @       @      @      &@                     �@@      U@       @      �?     �H@      (@     �w@      .@      f@      H@      @              �?      7@       @              ,@      "@     �X@      �?     �C@      $@      @              �?      ,@                       @              B@              9@      @      @                      "@       @              @      "@     �O@      �?      ,@      @                      @@     �N@              �?     �A@      @     �q@      ,@      a@      C@      �?              ;@      G@              �?      =@      �?     @m@       @     �W@      9@      �?              @      .@                      @       @     �G@      @     �E@      *@              ,@     @l@     @w@      :@      J@     v@     �P@     ��@     �g@     ��@     �m@      9@      @     �U@     @k@      &@      6@     @d@      >@     �w@      N@     Pt@     �[@       @      @     �K@     �Z@       @      $@     �V@      (@     �q@      D@     �i@     �Q@       @      @      B@     �I@      @      @     �O@      "@      W@     �A@     �V@      G@       @              3@      L@       @      @      <@      @      h@      @     @]@      9@                      ?@     �[@      @      (@     �Q@      2@     �X@      4@     �]@      D@      @              5@      I@       @      �?      @@      @      E@      @     @Q@      5@       @              $@     �N@      �?      &@     �C@      (@      L@      .@     �H@      3@      @      $@     �a@     @c@      .@      >@     �g@     �B@     `f@      `@     �i@     �_@      1@       @     �X@     @[@      (@      9@     �_@     �@@      U@     �X@      Z@     �U@      1@      @     �U@     @W@      &@      9@      \@      <@     �Q@     @R@      Y@      S@      @      �?      &@      0@      �?              ,@      @      *@      :@      @      &@      $@       @      E@     �F@      @      @     @P@      @     �W@      >@     �Y@     �C@                      0@      :@      @      �?      1@      @     �E@              8@      &@               @      :@      3@              @      H@      �?      J@      >@     �S@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ`�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?=��y@�	           ��@       	                    �?��>��d	@�           l�@                           �?��b:�@~           0�@                            �?[:��n@�            @o@������������������������       �Jt��@P            �_@������������������������       �:%=@�@G            �^@                            �?Fpt���@�            �v@������������������������       �탪��1@�            @m@������������������������       �-����@S            @`@
                           �?�����	@           ��@                            @ԓ\�;�	@�            �w@������������������������       �6�h9R	@q            `g@������������������������       �V��
�	@|            �g@                            �?ͩ�
�	@�           �@������������������������       �);U��
@�            �r@������������������������       �j�q3�@�            u@                          �4@�!�	@�           ܡ@                           �?!�]�h�@           $�@                          �0@��~�Ґ @-           �~@������������������������       �O@ o>_ @%            �P@������������������������       �MS��5 @           �z@                           @R��W�@�           ��@������������������������       ����o�@�             t@������������������������       �O�/C,@           �y@                          �7@V�D�ѱ@�           ��@                          �5@�#Qշx@V           ��@������������������������       ��*K�X@�            �i@������������������������       ��� 7�2@�            pt@                           @�$B�V@Q           ��@������������������������       �i$K�{�@!           |@������������������������       ����0@0            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@      t@     X�@      @@      I@     `|@     @V@      �@     �h@     �@     �x@     �@@      4@     �f@     �m@      9@      C@     `n@     �F@     �k@     �]@     �l@     �m@      8@       @     �I@     �V@      @      (@     �X@      &@      `@      B@     �W@     @T@      @      �?      7@     �G@       @      @     �M@       @     �E@      $@      <@      :@      @              "@      ?@               @      ?@      �?      2@      $@      ,@       @      @      �?      ,@      0@       @      @      <@      �?      9@              ,@      2@      �?      �?      <@     �E@      @      @     �C@      "@     @U@      :@     �P@     �K@       @      �?      *@      8@      @      @      6@      @     @P@      (@     �C@      E@                      .@      3@              �?      1@       @      4@      ,@      ;@      *@       @      2@     ``@     �b@      4@      :@      b@      A@     �W@     �T@      a@     �c@      2@      @      H@      N@      ,@      $@     �D@      0@      ?@      =@     �C@     @S@      @       @      :@      ?@      @      @      *@      (@      0@      2@      1@     �D@       @      @      6@      =@      &@      @      <@      @      .@      &@      6@      B@      @      *@     �T@     @V@      @      0@      Z@      2@      P@      K@     �X@      T@      (@       @      J@     �B@      @      "@      F@      $@      5@      <@      F@     �A@      @      @      ?@      J@      �?      @      N@       @     �E@      :@      K@     �F@      @       @     �a@     �s@      @      (@     `j@      F@     (�@     @S@     ؁@     �c@      "@             �N@      f@       @      @     �T@      @      @     �A@     �r@      O@      @              <@     �C@              �?      5@              n@      "@     �`@      1@      @                      $@                      @              <@              1@       @                      <@      =@              �?      1@             �j@      "@     �\@      "@      @             �@@      a@       @      @     �N@      @     �o@      :@     �d@     �F@                      3@     @R@      �?       @      C@      @     �T@      2@      N@      7@                      ,@      P@      �?      @      7@      �?     �e@       @     �Z@      6@               @     �S@     �a@      @      @      `@      D@     �n@      E@     q@     �W@      @             �B@      U@       @       @     @P@      8@     �b@      "@     ``@      <@       @              @      A@              �?      =@      .@      J@      @      L@      "@       @             �@@      I@       @      �?      B@      "@     @X@      @     �R@      3@               @      E@      L@      @      @      P@      0@      X@     �@@     �a@     �P@      @       @      9@      H@              @      K@      (@     �V@      ;@     �_@     �L@      @              1@       @      @              $@      @      @      @      0@      "@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @�~�$Q@�	           ��@       	                    �?11� 	@d           :�@                            �?A��YYj@�           ��@                          �;@��c@x            �g@������������������������       �f�]->D@j            �d@������������������������       ��3����@             ;@                          �<@l_�څ@.           �}@������������������������       �#1]b�@
            z@������������������������       ��&��N�@$             L@
                           @4�eQ�	@�           �@                           �?H�Ym�n	@F           0�@������������������������       ��˂rH�	@G            �[@������������������������       �1RJ�B;	@�           t�@                            @�`��	@x            @g@������������������������       ���$	@S            �`@������������������������       �l��Ѣ@%            �I@                           �?�_�@�@J           ��@                          �>@�(?`* @x            �@                           @?�fXh�?n           ��@������������������������       ��f|���?�            pw@������������������������       ���-O�y@{            �g@������������������������       ��:eϩ@
             .@                           @+�PF�@�           ��@                          �4@~�Qv��@�           �@������������������������       �
C�X��@a           X�@������������������������       �2�}�@]           Ȁ@                          �4@q� ѽ	@             B@������������������������       �fc��0�@             *@������������������������       �W=�{�@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        ,@     pq@     ��@      A@     �N@     �y@      V@     T�@     �n@      �@     �t@     �B@      (@      j@     0u@      ;@     �G@     �q@     �P@     `w@     �i@     �w@     �l@      ?@      @      N@     �V@       @      @     �O@      @     �d@     �C@     `d@      N@      @      @      ,@      A@              �?      .@       @      E@       @      N@      1@      �?              "@      ;@              �?      ,@      �?      E@       @      M@      $@              @      @      @                      �?      �?                       @      @      �?              G@     �L@       @      @      H@       @     @_@     �B@     �Y@     �E@      @              E@      J@       @       @     �C@       @     @^@      =@     @X@      9@      @              @      @               @      "@              @       @      @      2@              "@     �b@      o@      9@      E@     �k@     �O@     �i@     �d@      k@      e@      9@      @     �`@     �j@      8@     �D@      h@      H@     �g@     ``@     �i@     `c@      .@       @      $@      1@              (@      6@      @      @      (@      *@      &@      @      @     �^@     �h@      8@      =@     `e@     �F@     �f@     �]@     @h@      b@      &@       @      0@      A@      �?      �?      =@      .@      3@     �A@      $@      ,@      $@      �?      ,@      5@      �?              3@      .@      *@      :@      $@      @      "@      �?       @      *@              �?      $@              @      "@               @      �?       @     �Q@     �k@      @      ,@     @`@      5@     ��@     �D@     �z@      Y@      @              *@     �R@      �?      �?      :@      @      s@      &@      `@      *@       @              *@      R@      �?      �?      6@      @      s@      $@     �_@       @       @              "@     �F@                      ,@      @     �k@       @     @R@      @                      @      ;@      �?      �?       @             �T@       @      K@      @       @                       @                      @               @      �?      �?      @               @     �L@     �b@      @      *@      Z@      0@     �v@      >@     �r@     �U@      @       @      I@     @b@      @      $@      Y@      &@     �v@      :@     Pr@      U@      @              7@     �S@               @      D@      @      l@      (@     �a@      @@               @      ;@      Q@      @       @      N@       @      a@      ,@      c@      J@      @              @       @       @      @      @      @      @      @      @      @                              �?              @                      @              @      @                      @      �?       @              @      @              @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJlHachG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�2l@�	           ��@       	                    �?t���k�@W            �@                            �?��)8��@�           ��@                           �?��> u@�             w@������������������������       ����6�@�            0q@������������������������       ���P�d�@;            @W@                           �?�-"�E�@�            0r@������������������������       �ʁ���@W            @b@������������������������       ��y�,�@W             b@
                           �?~o�&	@�           ��@                          �5@�����	@�           x�@������������������������       �3Q�Jq�@0           0@������������������������       ��\��M/
@�           X�@                          �5@�D�c��@           �x@������������������������       �Q"�|@�             n@������������������������       �y�hdP@s            �c@                          �6@\.��@R           $�@                           �?��UT�@           �@                           �?�(Y�z�?'            ~@������������������������       �+�S���?�            0r@������������������������       �9&(�)�?            �g@                          �4@Q��ҧ�@�           ؆@������������������������       �i�E�&(@g           ��@������������������������       ��
E�@             i@                          �7@:�����@E           p�@                           @����@E            @]@������������������������       ��;@���@             E@������������������������       �o@-�j�@)            �R@                           �?�E��q@            �y@������������������������       �I�x��@@            �Z@������������������������       ���}Lr@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     `r@     x�@      @@     �O@      }@      Q@     ��@      m@     P�@     @v@     �@@      6@     `k@     �t@      6@      F@      t@     �J@     �u@     �g@     @v@     �n@      ;@      �?     �O@     �[@       @      &@     @T@      @      c@      9@     `a@     �N@      @      �?      =@     �M@              @     �@@      @     �V@      0@     �V@      A@      @      �?      8@      I@              @      =@      �?     �J@      ,@     @P@      =@      @              @      "@               @      @       @     �B@       @      :@      @      �?              A@      J@       @      @      H@      @      O@      "@      H@      ;@                      (@      9@       @      @      5@      @      ?@      @      8@      0@                      6@      ;@                      ;@              ?@      @      8@      &@              5@     �c@     @k@      4@     �@@     �m@      G@     �h@     �d@      k@      g@      5@      5@     @`@     �b@      .@      ;@     �f@     �B@     �\@     @^@     `c@     @b@      3@      "@      H@      L@       @      @     �T@      .@      R@     �G@     @W@     @P@       @      (@     �T@     �W@      *@      4@     �X@      6@     �E@     �R@      O@     @T@      1@              :@      Q@      @      @     �L@      "@     �T@      F@      O@      C@       @              @      G@      @      @      >@      @     @P@      ;@     �A@      4@                      5@      6@              @      ;@      @      1@      1@      ;@      2@       @       @     �R@     �l@      $@      3@      b@      .@     ��@      E@     `z@     �[@      @             �B@      c@      @      &@     @U@       @     p�@      0@     �r@      P@      @              (@      L@              @      6@      �?     p@      @     @\@      $@       @              @      =@              @      2@      �?     �d@      @      M@      @                      @      ;@                      @             �V@             �K@      @       @              9@     @X@      @      @     �O@      @     �p@      *@     @g@      K@      @              3@     @Q@      @      @     �A@       @      j@      *@     �`@      D@                      @      <@      @       @      <@      @      N@             �I@      ,@      @       @      C@     @S@      @       @     �M@      @     �`@      :@     �^@     �G@      �?              $@      @@              �?      @      @      B@      @      0@      @                      @       @                       @      @      (@       @      @       @                      @      8@              �?      @       @      8@      �?      $@      @               @      <@     �F@      @      @      J@       @     �X@      7@     �Z@      D@      �?                      $@                       @       @      C@      @      B@      @               @      <@     �A@      @      @      F@             �N@      1@     �Q@     �@@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��uk�C@�	           ��@       	                    �?.]��@}           H�@                           �?�<{�@@�           �@                           �?{R��@5           �|@������������������������       �R\���@}             h@������������������������       �rO�ԟ�@�            �p@                            �?��xCAH@m            �e@������������������������       ��� �@&             N@������������������������       �T�EO��@G            �\@
                           @)����y	@�           ��@                           �?4ы�;	@^           ��@������������������������       �>楍�y	@}           �@������������������������       �� T`�@�            �u@                           �?����`�	@}            �h@������������������������       �f@%�r�@            �J@������������������������       ��kѿ�@_            @b@                          �4@p��ǭ�@:           ��@                           �?^PO%�@G           8�@                          �0@����O�?�            `u@������������������������       �P>	�x�?!             K@������������������������       ��=���?�             r@                            �?3`n"@p           ��@������������������������       �f��q�&@�             w@������������������������       �^qY��@�            �k@                           �?-�!�~R@�           ��@                           �?�.��@�            @p@������������������������       �@ԢM�@]            @a@������������������������       �n�8f��@P            �^@                          �6@i�d$�@F           �@������������������������       �� �@x            �f@������������������������       �+ݫ��@�            Pt@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �q@     �~@      @@      J@     p@      S@     ؏@     �j@     �@     �u@      ?@      7@     �j@     �r@      8@     �E@     pu@     �N@     0x@     @e@     0w@     `o@      7@              L@     �T@       @      @     �S@      @     `e@     �A@     �a@      J@      @              D@     �Q@       @      @      L@      @     �[@      =@     �W@     �G@      @              4@      9@                      6@              M@       @     �D@      1@      �?              4@     �F@       @      @      A@      @      J@      5@     �J@      >@       @              0@      *@                      7@             �N@      @     �H@      @       @                       @                      @              2@              7@       @       @              0@      @                      0@             �E@      @      :@      @              7@     �c@     �k@      6@      B@     �p@     �L@      k@     �`@     �l@     �h@      2@      .@     �`@     @g@      4@     �A@     `m@     �F@     �g@     �Y@     `k@     �f@      *@      .@     �\@      `@      1@      ;@     �f@     �A@     @]@     �R@     �c@      b@      (@              4@     �L@      @       @     �J@      $@      R@      =@      N@     �B@      �?       @      6@      A@       @      �?      =@      (@      ;@      @@      "@      2@      @              (@      @                      ,@      @              @      @      "@      @       @      $@      ?@       @      �?      .@       @      ;@      <@      @      "@       @      @     @R@     �g@       @      "@      d@      .@     ��@     �F@     �|@      Y@       @              A@     @X@      @      "@     �M@      @     Pz@      4@     @n@      G@                      ,@      :@              @      &@              i@       @     �Q@       @                              $@                                      :@              0@       @                      ,@      0@              @      &@             �e@       @      K@      @                      4@     �Q@      @      @      H@      @     �k@      (@     �e@      C@                       @     �B@      @      @      C@             �a@      @     �\@      6@                      (@      A@      �?      �?      $@      @     @T@       @     �L@      0@              @     �C@     @W@      @             @Y@      (@     `j@      9@      k@      K@       @      @      "@     �B@                      6@       @     @X@      @     �P@      $@              @      @      3@                      1@      @      K@              A@      @                      @      2@                      @      @     �E@      @     �@@      @                      >@      L@      @             �S@      @     �\@      2@     �b@      F@       @              "@      5@      �?              6@      @      L@             �G@      *@       @              5@     �A@      @             �L@              M@      2@     �Y@      ?@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�}phG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �? �q��`@�	           ��@       	                    �?��XNMn@�           ��@                           �?5��R�@�           h�@                          �7@-篱�@�            �k@������������������������       �	)���@d            �b@������������������������       �6j4��X@/             R@                            �?��3� @           {@������������������������       �vI}w�>�?;            @Y@������������������������       �u31a�1@�            �t@
                          �=@�gQ�@X           ��@                           @����@L           8�@������������������������       ��A��-@�            ps@������������������������       ���Q�%� @�             j@������������������������       �W�3�-@             7@                           �?� B>�H@�           <�@                           @(aPYǪ	@�           �@                           �?�OKΊ	@�           ��@������������������������       ���J+F@�            �y@������������������������       ��� ���	@�           8�@                          �8@��aQ�@            �@@������������������������       �5"�$@             9@������������������������       �|R��>@              @                            �?�^�Y@�           h�@                           �?_�pWC�@�            Px@������������������������       �4�o��@h            `e@������������������������       ��ic�n@�            @k@                          �7@N��y}@�           T�@������������������������       �jK�'�@           Ȋ@������������������������       �$w.��@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        :@     �t@     ��@      =@      I@     �}@     �R@     ��@     �j@     Ї@     �w@      <@       @      Q@      d@       @       @     �[@      $@     �{@      C@     �p@     �T@      @       @      <@     �U@      �?      @      O@       @     q@      6@      _@     �D@      �?       @      1@      @@      �?      @     �D@      @      G@      *@     �A@      :@      �?              &@      6@                      <@       @      D@      "@      :@      "@      �?       @      @      $@      �?      @      *@      �?      @      @      "@      1@                      &@      K@               @      5@      @     `l@      "@     @V@      .@                              "@              �?      @      �?      O@              4@      @                      &@     �F@              �?      2@      @     �d@      "@     @Q@      $@                      D@     �R@      �?      @      H@       @     @e@      0@     �a@      E@      @              D@     �R@      �?      �?     �D@       @      e@      (@     `a@     �C@       @              B@      E@              �?      @@              Q@      "@      V@     �@@       @              @      @@      �?              "@       @      Y@      @     �I@      @                                               @      @               @      @       @      @      @      8@     Pp@     Pw@      ;@      E@     �v@      P@     ȁ@      f@     @     �r@      6@      6@     �a@      d@      1@      6@     �g@     �D@     �`@      Z@      b@      d@      1@      1@      a@      d@      1@      6@     �f@     �D@     �`@     �Y@     �a@      d@      *@      @      5@     �P@      @      "@     @S@       @     �P@     �@@      M@     �O@      @      *@     �\@     �W@      ,@      *@     �Y@     �@@     �P@     �Q@     �T@     @X@      "@      @      @      �?                      "@              �?      �?      @      �?      @      @      @                              @              �?              @              @                      �?                      @                      �?      �?      �?      �?       @     �]@     �j@      $@      4@      f@      7@     0{@      R@      v@      a@      @              C@     �I@              @      B@      @     �_@      3@     �Q@      C@                      3@      9@              �?      9@              F@      *@      :@      2@                      3@      :@               @      &@      @     �T@      @     �F@      4@               @      T@      d@      $@      1@     �a@      1@     @s@     �J@     �q@     �X@      @             �I@     �`@       @      &@     �R@      &@     �o@      ;@     �k@     �N@      @       @      =@      ;@       @      @     �P@      @      K@      :@     �N@     �B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��AhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?s�4��@�	           ��@       	                   �8@'�SW@�           4�@                          �2@cK��@k           ��@                            �?K�� @�            0y@������������������������       ����J� @z            �g@������������������������       �g�aW� @�            �j@                           �?���wD @l            �@������������������������       �(�/��@�             m@������������������������       ��-8#s@�            �u@
                          �<@C�s�T@�            �n@                          �9@�ݬ,io@X            �b@������������������������       ��'����@            �F@������������������������       ��c����@B             Z@                           �?��]3��@9            @X@������������������������       ��M�#�-@            �I@������������������������       ��g�ϟ@             G@                           @]p��@�           ��@                           @��NM	@�           ��@                           �?�\8��@M           ��@������������������������       ����N�
@L             ^@������������������������       �j/�T��@           �@                           �?(&�2��	@w            `e@������������������������       �(>#�[@!            �G@������������������������       ��pg	@V             _@                            �?�aaa��@�           P�@                           @�,q;@�            �@������������������������       ���_x�@�           ��@������������������������       �]<����@             (@                           �?JM絧�@H           ��@������������������������       �;��Zҙ@             B@������������������������       ��i����@3           �~@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@      �@      :@     �Q@     py@     �R@     ��@      h@     ��@      u@      =@      �?     @U@     �c@      @      (@     �U@      "@     }@     �B@     �q@     �S@      @             �P@      `@      @       @      J@      @     �y@      5@     �l@      I@      @              2@      ;@              @      ;@      �?     @j@      $@     @U@      6@                      &@      1@              �?      ,@             �W@       @      D@       @                      @      $@               @      *@      �?     �\@       @     �F@      ,@                     �H@     �Y@      @      @      9@      @     �i@      &@     �a@      <@      @              =@      F@      @      �?      *@             �G@      "@     �N@      3@      @              4@      M@      �?      @      (@      @     �c@       @     �T@      "@              �?      2@      >@              @     �A@      @     �I@      0@      L@      <@       @      �?      $@      4@                      8@      @     �A@      @     �E@      @       @              @      @                      @              &@      @      "@      @       @      �?      @      .@                      2@      @      8@       @      A@      �?                       @      $@              @      &@       @      0@      $@      *@      7@                      @       @              @               @      "@       @      @      1@                       @       @              �?      &@              @       @      "@      @              2@      k@     z@      3@      M@      t@     �P@     ��@     �c@     ��@     @p@      8@      *@     @c@      n@      *@     �E@      l@      K@     @l@      ^@     �k@     �f@      6@      $@     @a@      k@      (@      D@     �h@     �D@     �i@     �U@     `j@     �d@      *@      @      0@      "@              (@      5@      @      "@      &@      ,@      *@      @      @     �^@      j@      (@      <@     @f@     �A@     �h@      S@     �h@      c@       @      @      0@      7@      �?      @      :@      *@      3@     �@@      $@      .@      "@              @      @               @      (@      @      �?      @      @      @              @      "@      1@      �?      �?      ,@      "@      2@      =@      @       @      "@      @     �O@      f@      @      .@     �W@      (@     w@      B@     �s@     �S@       @             �B@     @W@       @      @      C@      @     �j@      7@      f@     �F@                     �B@     @W@      �?      @     �B@      @     �j@      6@     �e@     �E@                                      �?              �?      @              �?      @       @              @      :@      U@      @       @     �L@      @     @c@      *@      a@      A@       @      @      @      "@              �?      @      @       @      @      @                              7@     �R@      @      @      K@       @      c@      "@     @`@      A@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���^hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�a�^@�	           ��@       	                    @�u�\ͬ@q           ��@                          �2@h.��@�           ܐ@                           �?��nh{C@+           `|@������������������������       ��R��@�            `t@������������������������       ��yL�@Z             `@                          �4@��5Нw@�           ��@������������������������       �P��@�@            z@������������������������       ��V�[χ@�            �i@
                           @u"\u@�           ��@                           @�_s"��@�            `p@������������������������       �-U�k�Q@�            `j@������������������������       ��O (Y�@             �I@                            �?�^�8�@           Ј@������������������������       ��	��~:�?j            �c@������������������������       ���I@�           ��@                           �?�g	b��@d           ț@                            �?����@%           @|@                           �?�&��"�@Q            �^@������������������������       ���?��\@#            �J@������������������������       ��s���@.            @Q@                          �@@���$�@�            �t@������������������������       �jv� w@�            �s@������������������������       ���^~@             &@                           @���S	@?           ��@                           �?ܮ_��	@           ��@������������������������       �[ji�@/             R@������������������������       �/Aq��	@�           @�@                           @2`�@4           �}@������������������������       �#s�wYS@*           �|@������������������������       �`2s?��?
             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@      s@     x�@      <@      P@     P{@     �V@     ��@     �k@     `�@     �v@     �@@      @     @_@      s@       @      B@      i@     �C@     ��@      V@     @|@     �b@      "@      @     �T@     �d@      @      5@     @a@      ;@     @o@      S@      i@     @Y@      @       @      A@     �P@              @     �P@      @     �_@      7@     @T@     �F@               @      =@     �H@              @     �J@      @     @R@      .@     �M@      B@                      @      1@              �?      *@             �J@       @      6@      "@              @      H@     @Y@      @      .@      R@      6@      _@     �J@      ^@      L@      @       @      <@      L@      @       @     �I@      .@     �V@      C@      S@      E@      @      �?      4@     �F@              @      5@      @     �@@      .@      F@      ,@                     �E@      a@      @      .@     �O@      (@     `}@      (@     `o@     �G@      @              1@     �H@                      .@      &@     �V@      @     �N@      .@      �?              $@      D@                      .@      "@     �Q@              J@      ,@                      @      "@                               @      3@      @      "@      �?      �?              :@      V@      @      .@      H@      �?     �w@      "@     �g@      @@       @               @      $@              @      &@             �W@              >@       @                      8@     �S@      @      (@     �B@      �?     �q@      "@      d@      8@       @       @     `f@     �o@      4@      <@     �m@      J@     �r@     �`@     �t@     �j@      8@      �?      C@     �P@              @     �J@      @     �[@      0@     �]@      D@      �?      �?      (@      8@               @      2@      @      6@      @      >@      @      �?      �?      @      @               @      @       @      .@       @      "@      @                      @      1@                      &@      �?      @      �?      5@      @      �?              :@      E@               @     �A@      �?     @V@      *@      V@      A@                      :@      E@                      ?@      �?     @V@      &@     �U@      @@                                               @      @                       @      �?       @              @     �a@     �g@      4@      8@     �f@      H@     �g@     @]@     @j@     �e@      7@      @     �V@     �a@      .@      3@     �\@      C@     @R@      Y@     �X@     @`@      6@       @      &@      *@              @      1@      @              $@      @      @      �?      @      T@     �_@      .@      *@     �X@     �A@     @R@     �V@     @W@     �_@      5@      �?      I@     �H@      @      @      Q@      $@     �]@      1@     �[@     �E@      �?      �?     �D@     �H@       @      @     @P@      $@     @]@      ,@     �[@     �E@      �?              "@              @              @              �?      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�)�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�G�@,@@�	           ��@       	                    �?��pu��@�           h�@                           �?�y��H@�             t@                          �<@r��@̹@e            �c@������������������������       ����+x@\            �a@������������������������       �i	\��p @	             0@                          �4@n�U%�@o            �d@������������������������       ��f?iun�?<            @W@������������������������       ��{�N��@3             R@
                           �?�2��1�@�           X�@                          �:@�V	@�            �r@������������������������       � ���@�            @l@������������������������       ��\�W��@-            @R@                          �5@U@Ii@�             x@������������������������       �6�/���@�             k@������������������������       ��rlz@e            �d@                          �5@��hW�b@           ��@                          �1@�;�xF�@�           <�@                           @S�d���@           �z@������������������������       �YE���B@q            �d@������������������������       ����s��?�            0p@                            �?ò��!�@�           ��@������������������������       ��
��X�@'           �}@������������������������       ��ll�/@�           H�@                           @�"��,�@           4�@                           @��D�Q_@�           �@������������������������       �Gu�J�O	@�           ��@������������������������       �%e^a�V@           �z@                          �;@A�hb��@R             b@������������������������       �
g� ��@?             Y@������������������������       �7��[C:@            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pq@     h�@      8@      L@     p~@     @U@     ��@      k@     x�@     �t@      <@       @     �T@     �`@      @      &@     �\@      0@     �r@     �L@     `g@     @V@      "@              ,@     �G@               @      8@      @     �`@       @      Q@      2@      �?              @      2@               @      .@      @      S@      @      9@      @                       @      (@               @      .@      @      S@      @      4@      @                       @      @                              �?                      @       @                      $@      =@                      "@      �?     �M@       @     �E@      &@      �?              @      $@                      �?             �G@      �?      7@      @                      @      3@                       @      �?      (@      �?      4@      @      �?       @     @Q@     �U@      @      "@     �V@      &@     `d@     �H@     �]@     �Q@       @       @      C@     �C@      @      @     �I@      @     �C@      A@     �E@      <@       @      �?      B@      ?@      @      @     �C@       @      =@      3@      B@      3@      @      �?       @       @              @      (@      @      $@      .@      @      "@      �?              ?@      H@       @       @     �C@      @      _@      .@      S@     �E@                      @      ?@              �?      3@             @T@      @      K@      6@                      ;@      1@       @      �?      4@      @     �E@      $@      6@      5@              4@     �h@     p|@      3@     �F@     Pw@     @Q@     0�@      d@     ��@     �n@      3@       @      T@     �n@      "@      .@     �d@      @@     �@     �Q@     `v@      ]@      @       @      4@     @P@      �?      �?     �A@             `f@      (@      V@      5@      �?       @      0@      <@      �?      �?      4@              H@      (@      9@      *@                      @     �B@                      .@             ``@             �O@       @      �?      @      N@     �f@       @      ,@     ``@      @@     �t@      M@     �p@     �W@      @       @      =@      W@      @      @     �F@      &@     @[@      3@     �]@      A@      @      @      ?@     �V@      �?       @     �U@      5@     `k@     �C@     �b@     �N@       @      (@      ]@      j@      $@      >@     �i@     �B@     `i@     �V@     �m@     @`@      (@      @     �Y@     �f@      "@      >@      f@     �A@      g@     �O@     �l@      _@       @      @      T@      ^@      @      :@     @]@      @@     �V@     �H@     �X@     �V@       @      �?      7@      O@      @      @     �M@      @     �W@      ,@      `@      A@              @      *@      :@      �?              ?@       @      3@      ;@      $@      @      @       @       @      2@      �?              $@       @      3@      8@       @      @      @      @      @       @                      5@                      @       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Di4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@| o�_X@�	           ��@       	                    �?��ti@P           ��@                           �?��O��@�           ��@                            �?:p��@�            �p@������������������������       �O��@,            @P@������������������������       �~�-�@�            �i@                           �??��@<           p~@������������������������       �#�V^Ó@l             e@������������������������       �#���^{@�            �s@
                           @�pL�
?@h           $�@                          �0@�ʖ�[i@�            Pv@������������������������       ���uw�� @             C@������������������������       �f���@�            �s@                          �4@?��J�@�           ��@������������������������       ��W�ǁ)@5           ��@������������������������       ��}`Â�@_             e@                          �<@�-JH�@E           (�@                          �9@a���@w           �@                           �?%�p�a@y            �@������������������������       �����w	@           �{@������������������������       ������@Z           (�@                           �?���qM�@�            �y@������������������������       ��E�	@�            �j@������������������������       �0E����@~            `i@                            �?�� 	@�            pt@                           @��Ix*@n            �e@������������������������       ��h��P�@D            @Z@������������������������       �]B�'G�@*            �Q@                           �?��{���@`             c@������������������������       �,M#�@#            �H@������������������������       �	^Δo@=            �Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �r@     ��@     �@@     �H@     }@     @S@     ��@     �l@     ��@     pv@      =@      (@     @]@     @r@      "@      3@     �h@      3@     ؅@     @[@     ��@     `d@      "@      (@      O@     @V@      @      $@     @Y@      $@     �d@     �Q@     �a@     �U@      @              .@     �E@      �?       @      8@       @     @S@      3@      N@      :@       @              �?      &@                      @              2@      �?      8@      @                      ,@      @@      �?       @      4@       @     �M@      2@      B@      4@       @      (@     �G@      G@      @       @     @S@       @     �V@      J@     @T@      N@       @      @      ,@      3@      @      �?      ?@      @      <@      .@      ;@      5@              @     �@@      ;@      �?      @      G@      @      O@     �B@      K@     �C@       @             �K@     `i@      @      "@     �X@      "@     ��@      C@     0x@     @S@      @              .@     @P@      �?       @      A@      �?     �[@      6@     �U@      4@                      �?      0@                      @              @              "@      �?                      ,@     �H@      �?       @      >@      �?      Z@      6@     @S@      3@                      D@     @a@      @      @      P@       @     Pz@      0@     �r@     �L@      @              C@     �Y@      @      @      K@       @      w@      ,@     `o@     �I@      �?               @     �A@               @      $@      @     �I@       @      I@      @      @      *@     �f@      n@      8@      >@     �p@      M@     0r@     �]@     �r@     �h@      4@      @      b@     �g@      2@      :@     �i@      E@     �p@     �V@     �p@      a@      2@      @      ]@     �a@      "@      6@      c@      9@     �f@     �J@     �f@     @X@      *@       @      O@      Q@      @      ,@     @S@      *@      D@     �C@     @Q@      F@      (@      �?      K@     �R@       @       @     �R@      (@     �a@      ,@      \@     �J@      �?      @      <@      H@      "@      @     �K@      1@     �T@      C@      U@      D@      @      @      *@     �@@      @      �?      =@      1@      <@      3@     �@@      8@      @              .@      .@      @      @      :@             �K@      3@     �I@      0@              @     �B@      I@      @      @     �M@      0@      9@      <@     �A@     �M@       @      �?      (@      4@               @      ;@      &@      (@      5@      8@     �E@       @              @      ,@               @      1@      $@      @      $@      @     �A@       @      �?       @      @                      $@      �?      @      &@      3@       @              @      9@      >@      @       @      @@      @      *@      @      &@      0@              @      @      ,@       @       @      $@      �?      @      �?      @      @                      6@      0@      @              6@      @      $@      @       @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�W�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�c�d>@�	           ��@       	                    �?b��Y�@{           N�@                           �?�p����@           ��@                           @�ܿٔ@�            Pp@������������������������       �J��"�@�            �l@������������������������       ���p`�@             >@                          �;@ukr	@           x�@������������������������       ���/n�@H           0@������������������������       �ܝ9��@7             W@
                           �?l���Di@^           L�@                           �?�&�`I�@�            �t@������������������������       ���᧿o@�            @n@������������������������       �aN�y�@:            @W@                           �?����	@�           �@������������������������       � OM;% @=            �U@������������������������       �zf&b)�@I           h�@                          �1@ �M.@1           ��@                           @��8$ @�            Pv@                           @T�n!��?�            @q@������������������������       �}����?T            �`@������������������������       ��jH�7j�?X            �a@                           �?\�V�L@-            @T@������������������������       �
.�x��@             D@������������������������       �'F<7VZ@            �D@                          �5@�T��s�@X           ��@                           @�񳴙@�           X�@������������������������       �#�鰂@u            �h@������������������������       �����x@e           (�@                          �8@:�D@~           ��@������������������������       �ϋ�Zݸ@�            �r@������������������������       ���hí@�            Pr@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      r@     ��@      <@      F@     �|@     @W@     Ў@     `k@     `�@     @u@      ?@      2@      h@     �u@      2@     �A@     �s@     @Q@     pw@      f@     �x@     �n@      9@      @      R@     �c@      &@      ,@      _@      ;@     �b@     �M@     �^@     �W@      .@       @      ,@     �G@       @      @      L@       @     �J@      @      C@      9@      @       @      "@     �G@       @      @      F@       @     �J@      @     �B@      6@      @              @                              (@      @              �?      �?      @       @      @      M@     �[@      "@      $@      Q@      3@     @X@      K@      U@     @Q@       @      @      K@     �W@      "@      "@      H@      *@     �V@     �E@     �S@      I@       @       @      @      0@              �?      4@      @      @      &@      @      3@              &@      ^@     �g@      @      5@     `h@      E@      l@     �]@      q@     �b@      $@             �E@     �D@                     �C@              T@      "@     �W@      <@      �?             �A@      B@                      A@              J@       @      K@      6@      �?               @      @                      @              <@      �?      D@      @              &@     @S@     �b@      @      5@     �c@      E@      b@     @[@     �f@     �^@      "@      @      $@      @              @      1@      �?      @      $@      3@      (@              @     �P@      b@      @      .@     `a@     �D@     �a@     �X@      d@     �[@      "@       @     �X@     �j@      $@      "@     @a@      8@     �@      E@      |@     �W@      @              @     �@@               @      6@              h@      @     @S@      1@      @              @      9@                       @             �d@      �?      L@      ,@                      @      *@                      �?             �W@              3@      @                      �?      (@                      @             @R@      �?     �B@      &@                      �?       @               @      ,@              :@      @      5@      @      @                      @               @      $@              .@              @      @                      �?      @                      @              &@      @      ,@              @       @      W@     �f@      $@      @      ]@      8@      z@      C@     0w@     �S@      @              G@     �[@       @      @     �G@      .@     �p@      2@     @j@      :@       @              <@     �D@                      .@      @      G@      $@     �D@       @       @              2@     �Q@       @      @      @@       @     �k@       @      e@      2@               @      G@     �Q@       @      @     @Q@      "@      c@      4@      d@      J@      �?       @      =@      B@      @      �?     �B@      @     �W@      @     �O@      :@      �?              1@     �A@      @       @      @@      @      M@      1@     �X@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?ӓ�
]=@�	           ��@                           �?���;&�@           h�@                           @@~�ls'@2           p@                          �;@H���@)           P~@������������������������       ��m�Q?@           �z@������������������������       �H����	@#             M@������������������������       �6�:����?	             2@                           @�%�r��@�           �@	       
                   �4@�l�,��@�             r@������������������������       �`kt� @g             b@������������������������       �>G4�L�@[            @b@                            @���c3� @           |@������������������������       �m�X@�            @w@������������������������       �1�&J��?2            @S@                           @NpD�@�           ޤ@                           �?$��7	@�           t�@                           @	+�*�	@�           ��@������������������������       ��3�o	@|           H�@������������������������       ����a	@W            @_@                           �?B��"�@           p{@������������������������       ��7�8q#@j            `d@������������������������       ��z ڼ@�            @q@                          �7@B�r^�@�           H�@                          �6@Z/K�P�@           ��@������������������������       ��~j��@@�           p�@������������������������       �|���@.            �Q@                            @���7�e@�            �q@������������������������       ��[>xFe@�            �k@������������������������       �ݺ�B{@%             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        .@     �r@     ��@      4@      K@      }@     �W@     ��@      l@     ��@     �v@      9@      @     �Q@     �e@       @      .@     �Z@      0@     �{@      E@     @r@     @S@      @      @     �C@     �T@      �?      *@     @R@      @     �\@      ;@     �X@     �G@      @      @      C@      T@      �?      @     �P@      @     �\@      ;@      X@     �G@      @             �A@      R@      �?      @      O@       @     @Z@      7@     �U@     �@@      @      @      @       @               @      @      �?      "@      @      "@      ,@                      �?       @              @      @                               @                              ?@     �V@      �?       @      A@      *@     �t@      .@     @h@      >@      �?              1@      A@                      ,@      (@     �]@      @     �R@      0@      �?              &@      ,@                      @             �P@      �?      E@      @                      @      4@                      $@      (@     �I@       @     �@@      &@      �?              ,@      L@      �?       @      4@      �?     @j@      (@     �]@      ,@                      (@     �K@      �?              1@      �?     @d@      &@      Y@      *@                       @      �?               @      @              H@      �?      3@      �?              (@      m@     0w@      2@     �C@     pv@     �S@      �@     �f@     h�@     �q@      5@      (@     `d@     �m@      *@      A@     �m@     �O@     @h@     �c@     �m@     �h@      1@      (@     �_@      d@      (@      ;@      f@      H@      ]@     �]@     �c@     @c@      1@      "@     �[@     �a@      &@      ;@     @c@      E@     �Y@      X@      c@     �a@      &@      @      .@      1@      �?              7@      @      *@      7@      @      *@      @             �B@     �S@      �?      @     �N@      .@     �S@      D@      T@      E@                      &@      ;@               @      6@      @      :@      2@     �A@      2@                      :@     �I@      �?      @     �C@      &@      J@      6@     �F@      8@                     �Q@     �`@      @      @     @^@      .@      v@      7@     �q@     @V@      @             �C@     �Z@      @      @      P@      $@      s@      &@     �k@      K@      @              A@     �U@      @      @     �M@      @      r@      &@      i@      J@      @              @      4@              �?      @      @      ,@              3@       @                      ?@      :@       @             �L@      @      I@      (@     �P@     �A@      �?              >@      6@                     �E@      @     �A@      "@      I@      ;@      �?              �?      @       @              ,@              .@      @      1@       @        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @��2�w�@�	           ��@       	                   �<@G�n@j	@�           ��@                          �2@kH@�@�           �@                           @��L��g@+           �|@������������������������       �C(o�F�@           �z@������������������������       �s4Y�m@             ?@                           �?/oHz�(	@�           ��@������������������������       �zXբ	@�           P�@������������������������       �sш� +@�            �y@
                          �A@m�e)�	@�            `q@                          �?@U���"�	@�             p@������������������������       ��
�7	@p            �g@������������������������       �]o�}@+            �P@������������������������       ����G��@
             4@                           �?1du:�M@           �@                           @��Kڣ� @U           �@                           @�[�5E�?�            pr@������������������������       �18���@W             a@������������������������       �zR[���?c            �c@                           �?�c�)!N@�            `o@������������������������       �L{?�m�@[             b@������������������������       �?Q����?@            �Z@                          �7@J�2�~@�           `�@                           �?>�%S�@           ��@������������������������       �k�!u�@�            `y@������������������������       �s�����@
           z@                            �?Q�t�@�            r@������������������������       ����H@V            �`@������������������������       ���Ö:@\            @c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        5@     �s@     ��@      A@     �K@      ~@     �X@     ؍@     �k@     x�@     �w@      A@      5@      l@      s@      :@      D@     pt@     �S@     v@      h@     �x@     �p@      =@      (@      i@      q@      8@      ;@     `r@     �M@     �u@      c@     Pv@      j@      8@      �?      C@      O@              @      O@      @      \@      @@      W@      K@      �?      �?     �A@      N@              @     �J@             �[@      <@     @V@      I@                      @       @                      "@      @       @      @      @      @      �?      &@     `d@     �j@      8@      8@      m@      L@      m@      ^@     �p@     `c@      7@      &@     @`@     �b@      7@      2@     �e@      F@     �b@     @W@     �f@      ]@      7@             �@@      P@      �?      @      N@      (@     �T@      ;@      U@     �C@              "@      8@      @@       @      *@     �@@      3@      "@      D@      B@      L@      @      @      8@      9@       @      *@      ?@      3@      "@     �C@      A@     �J@      @       @      (@      6@              &@      3@      *@      "@      <@      =@     �D@      @       @      (@      @       @       @      (@      @              &@      @      (@              @              @                       @                      �?       @      @                      V@     �l@       @      .@     `c@      5@     Ђ@      ?@     `x@     �\@      @              (@     �P@              @     �A@       @     `q@      @     @^@      0@       @               @      A@                      (@       @     �d@      @     �K@       @                      @      5@                      "@      @     �N@       @      =@      @                      @      *@                      @      @     �Z@      �?      :@      @                      @      @@              @      7@             �[@       @     �P@       @       @              @      6@              @      (@             @Q@       @      <@      @                              $@                      &@              E@              C@      @       @              S@     @d@       @      (@      ^@      *@     @t@      :@     �p@     �X@      @              J@     @`@      @      @      T@      $@     �p@      *@     �i@     �I@      @              ?@      M@      �?      @      N@       @     �]@      @     @Y@      5@      @              5@      R@      @       @      4@       @     �b@      @      Z@      >@                      8@      @@      @      @      D@      @     �L@      *@      P@      H@                       @      2@               @      "@              :@       @     �A@      =@                      0@      ,@      @      @      ?@      @      ?@      @      =@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ6aKhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�PE�yP@�	           ��@       	                   �3@X�`��@L           ��@                           �?2)P�@�           ��@                          �1@�}��^@�             o@������������������������       ��{��@<            @X@������������������������       ����@b             c@                          �1@I�60@           �{@������������������������       �oG2_�z@j            `e@������������������������       �~����@�             q@
                           �?8�b)	@�           \�@                          �<@����@�            Px@������������������������       ��{�y�@�            �t@������������������������       �*jg���@'             K@                           @u�&Л�	@�           H�@������������������������       �-a�n|�	@=           ��@������������������������       ���A;)�	@\            �c@                           @u��@Z           ��@                          �1@kp��)@           �y@                            �?��1�.��?6             T@������������������������       �X��Ce�?             :@������������������������       �r���W_�?%             K@                          �7@|��(�@�            �t@������������������������       ���C��^@�            `l@������������������������       ��h���@B             Z@                          �5@h�E t�@S           ��@                           @V<�&ܵ@"           ��@������������������������       ���	W @V           0�@������������������������       ���D�@�            �t@                           @s���@1            @������������������������       �"���@�            `o@������������������������       ��ʑ��@�            �n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �p@     ��@     �F@     �E@     �{@     �U@     �@      j@     (�@     �v@     �@@      6@     �f@     �t@     �@@      >@     �r@      O@     �v@      f@     0v@     �m@      ;@      @     �D@     �W@      @      @     @U@      2@     `f@      I@     @`@      T@       @              &@      A@                      ;@      @     �T@      "@     �M@      5@                      @      (@                      (@             �E@      @      3@      @                       @      6@                      .@      @      D@      @      D@      2@              @      >@     �N@      @      @      M@      *@      X@     �D@     �Q@     �M@       @      �?      &@      >@      �?       @      $@       @      G@      ,@      @@      6@              @      3@      ?@       @       @      H@      &@      I@      ;@     �C@     �B@       @      1@     �a@     �m@      >@      :@      k@      F@      g@     �_@      l@     �c@      9@      �?     �A@      O@      �?      @      I@      @     �U@      :@     �T@      A@      @      �?     �@@     �I@      �?      �?      D@      @     �T@      3@     @S@      4@      @               @      &@               @      $@              @      @      @      ,@              0@     @Z@     �e@      =@      7@     �d@      C@     �X@     @Y@     �a@      _@      6@      @     �U@     �b@      :@      6@     �b@      @@     �T@     @Q@     �`@     @[@      3@      $@      3@      8@      @      �?      2@      @      1@      @@       @      .@      @       @      V@     @m@      (@      *@     �a@      9@     ��@      ?@      |@     �^@      @       @      A@     @Q@      �?              @@      0@     �`@      @     �U@      @@       @               @       @                      �?              G@      �?      1@      @                                                                      3@      �?      �?      @                       @       @                      �?              ;@              0@                       @      @@     �N@      �?              ?@      0@     �U@      @     @Q@      ;@       @              5@     �I@      �?              ,@      *@     �P@       @      D@      0@       @       @      &@      $@                      1@      @      4@      �?      =@      &@                      K@     �d@      &@      *@     �[@      "@     ��@      ;@     �v@     �V@      @              8@     �V@      @      $@      L@       @     �x@       @     �m@     �G@      @              ,@     �K@       @      @      <@             �p@      @     �c@      3@                      $@     �A@      @      @      <@       @     �`@      @     @T@      <@      @              >@     �R@      @      @      K@      @     �`@      3@     �_@      F@      �?              0@      C@              �?      6@             @U@      @      O@      3@      �?              ,@     �B@      @       @      @@      @     �G@      (@      P@      9@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�/XhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�$��o@�	           ��@       	                    �?��o!`	@           ��@                           �?G *`�@6           ~@                            @_�qF@~            `g@������������������������       �2���@\             a@������������������������       �>n�6\:�?"             I@                           �?da9�@�            `r@������������������������       �
���id	@W            �b@������������������������       �6L8��@a             b@
                          �:@��#V�	@�            �@                           �?��~|�	@A           (�@������������������������       � �ནn	@�            �t@������������������������       �gC��l	@}           ��@                           �?��G�C�@�            `o@������������������������       �a>:|�@.             R@������������������������       �$mWl@u            `f@                           @X����@�           С@                            @�c<�@l           ȁ@                          �3@�2�6<+@
           0z@������������������������       �t{!�<�@d            `d@������������������������       �"�(_�@�             p@                           �?��-nS@b            �b@������������������������       ��ң45�?             A@������������������������       �!O<q@I             ]@                          �6@ަ��$@D           ��@                           �?��v�tY@           ��@������������������������       �?����@�           ��@������������������������       ��'8�(�@i           ��@                          �<@�H��`�@B           �@������������������������       ���@           @z@������������������������       �ܫ� W@<            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     (�@      @@     �J@     �{@     �R@     �@      m@      �@     �x@     �@@      0@      f@     �n@      4@     �@@     �m@     �H@     �j@     `a@      o@     �k@      ?@       @     �J@     @Q@       @      @      M@      @     �Y@      3@     �X@     �K@       @       @      .@      5@                      1@             �K@       @     �K@      2@       @       @      "@      .@                      0@             �@@       @      D@      2@       @              @      @                      �?              6@              .@                              C@      H@       @      @     �D@      @      H@      1@      F@     �B@      @              1@      4@       @      @      5@      @      9@      $@      1@      6@      @              5@      <@               @      4@              7@      @      ;@      .@       @      ,@     �^@      f@      2@      ;@     �f@      E@     �[@      ^@     �b@      e@      7@      @     �W@     @b@      &@      8@     �b@      B@     @W@     @W@      _@     @Y@      7@       @     �B@      S@      @      @      H@      *@      >@      @@      <@      C@      (@      @      M@     �Q@      @      2@     @Y@      7@     �O@     �N@      X@     �O@      &@       @      <@      ?@      @      @      ?@      @      2@      ;@      9@     �P@              �?      @      @       @      �?      $@              $@      &@      $@      4@              @      9@      ;@      @       @      5@      @       @      0@      .@     �G@                     �a@     �r@      (@      4@     �i@      :@     h�@     �W@     @�@     �e@       @              K@     �S@      @      "@     �N@      (@      b@     �F@      [@      K@                     �F@     �G@      �?       @     �J@      $@     @W@     �A@      W@     �A@                      .@      2@                      ,@              D@      .@     �G@      ,@                      >@      =@      �?       @     �C@      $@     �J@      4@     �F@      5@                      "@      ?@       @      �?       @       @      J@      $@      0@      3@                               @                      @              .@      �?      &@      �?                      "@      =@       @      �?      @       @     �B@      "@      @      2@                     @V@      l@      "@      &@      b@      ,@     ��@     �H@     �y@      ^@       @             �G@     @c@      @      @     �U@      "@     ��@      4@     �q@      M@      �?              7@     @R@       @      @      K@      @     �r@      @      `@     �A@      �?              8@     @T@      @             �@@      @     @l@      0@      c@      7@                      E@     �Q@      @      @     �L@      @     �Z@      =@     �`@      O@      �?              >@      L@      �?      @      @@      @      X@      =@     �]@      I@      �?              (@      .@      @       @      9@      �?      &@              ,@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�N�'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�����P@	           ��@       	                   �;@2��+	@�           ��@                           �?�c��@L           ��@                          �1@R|:��@K           ��@������������������������       ��/_R<I@7            �U@������������������������       ���v�O@           �{@                           @��R2�J	@           h�@������������������������       �X��+�@;           h�@������������������������       ��͕�lt	@�             t@
                          @@@L�%y	@�            �p@                            �?�}��$	@�            �j@������������������������       ��"�a��	@%             I@������������������������       ��o���@h            `d@                            �?W�(���@            �K@������������������������       �i�T���?             1@������������������������       �|����!@             C@                           @�}Q���@�           ��@                          �7@��$���@h           �@                           @ˁKLM�@�            `y@������������������������       ��n��K�@l             e@������������������������       ��ĉ�W@�            �m@                            @�����@m            �e@������������������������       ��V	J;Q@E            �[@������������������������       �:�t�'�@(            �N@                            �?��(@!           h�@                            �?̽�4�/@A           ��@������������������������       �`rd�@�            �x@������������������������       ��O��i@Q           `�@                           �?�����@�           �@������������������������       ����D�h@�            �p@������������������������       �U�cE�@4           P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      q@     @�@      >@      Q@      |@     @R@     ��@     �k@     H�@     �w@      4@      6@     `d@     �m@      5@     �E@     �n@      F@      k@      a@     �q@     `k@      *@      $@     `a@     �h@      2@      B@      j@     �A@     �h@     @]@     �o@      c@      &@      �?     �B@     �T@       @      *@     @R@      &@     �W@      D@     �Z@     �P@      @              @      @                      @      �?      <@       @      7@      $@              �?      A@     �R@       @      *@     �P@      $@     �P@      @@      U@      L@      @      "@     �Y@     �\@      0@      7@      a@      8@     �Y@     @S@     �b@     �U@      @      �?      Q@      R@      ,@      1@     �U@      .@      R@      B@      Y@     �E@      �?       @      A@      E@       @      @      I@      "@      ?@     �D@      H@      F@      @      (@      8@      D@      @      @     �A@      "@      3@      3@      @@     �P@       @      @      3@      =@      @      @      <@      @      3@      3@      5@      K@       @              �?       @      �?      @       @      @      @       @      @      @       @      @      2@      5@       @      @      4@       @      *@      &@      1@     �H@              @      @      &@              �?      @      @                      &@      (@                              @                      @                                      @              @      @      @              �?      @      @                      &@      @              �?     �[@     �u@      "@      9@     �i@      =@     ؇@     �U@     P�@     @d@      @              A@      W@      �?      $@     @S@      "@      c@     �E@      Z@      K@       @              4@     �O@      �?       @     �N@      @     @^@      4@     �S@      =@      �?              &@      0@              @      >@             �P@       @      <@      (@                      "@     �G@      �?      @      ?@      @     �K@      2@     �I@      1@      �?              ,@      =@               @      0@      @      ?@      7@      9@      9@      �?              @      ,@               @      *@      @      .@      2@      2@      1@      �?              @      .@                      @              0@      @      @       @              �?     @S@      p@       @      .@     �_@      4@     �@      F@      z@      [@      @              E@     @a@      @      *@     @P@      (@     @t@      8@      m@     �P@                      1@     �J@       @      @      8@      @     `d@       @     �T@     �B@                      9@     @U@      �?      $@     �D@      @      d@      0@     �b@      >@              �?     �A@     �]@      @       @      O@       @     �q@      4@     @g@     �D@      @      �?       @      E@                      (@      @     �^@      ,@      P@      @                      ;@      S@      @       @      I@      @     �d@      @     �^@      C@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��uthG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�%��\@�	           ��@       	                   �8@�/C�@�           T�@                           �?�����@�           h�@                           �?L�C�@7           ~@������������������������       �&�L�,�@�            `v@������������������������       � �K�r@U            �^@                          �4@WI��7�@�           �@������������������������       ��~��!�@�           0�@������������������������       �X��:��@-           0}@
                           �?�D��$

@�           ��@                          �:@�8a�aA
@L            �@������������������������       ����M�@r            �e@������������������������       ������5
@�            @u@                            �?�3k�@U             b@������������������������       �X>sF�@             D@������������������������       �d�,7Ys@=             Z@                           �?�sn�@6           |�@                            @'�X";@e           �@                          �4@�2�u{�@3           �~@������������������������       ���V�L(�?�            @s@������������������������       �V�����@z            `g@                          �2@j� �v��?2             U@������������������������       �z#����?            �D@������������������������       �и:��+�?            �E@                          �7@�BR�y@�           p�@                           @(/��	�@           H�@������������������������       �����k�@Z           ��@������������������������       ��Eq㸔@�            @q@                           @������@�            0s@������������������������       ��=��@"             L@������������������������       �@0(�@�            `o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     pr@     �@      ?@      I@     P}@     �U@     h�@     @l@     Љ@     �v@      <@      2@     �j@     0s@      9@      D@     0t@     @Q@     �w@      g@     @x@      o@      9@      @     �_@     �k@      .@      :@      k@     �C@     �s@     �]@      s@     �d@      "@              =@     �P@      �?      @     �K@       @      `@      2@      `@      H@                      6@      L@      �?      @     �E@      �?     @T@      0@      W@     �E@                      @      $@              �?      (@      �?      H@       @     �B@      @              @     �X@     �c@      ,@      6@     @d@     �B@      g@      Y@     �e@      ]@      "@      @      H@     �Q@      $@       @     �V@      .@     @^@     �P@     @[@     @P@      @      �?      I@     �U@      @      ,@      R@      6@     �O@      A@     �P@     �I@      @      &@     �U@      U@      $@      ,@     �Z@      >@     �O@     �P@      U@     @U@      0@      &@     �K@     �N@      $@      *@     �V@      6@     �F@      L@     @P@     �Q@      ,@              7@      ?@       @      �?      =@      @      0@      9@      3@      &@      "@      &@      @@      >@       @      (@     �N@      0@      =@      ?@      G@     �M@      @              ?@      7@              �?      0@       @      2@      &@      3@      .@       @              @      $@                      @      �?      @               @      @       @              ;@      *@              �?      $@      @      ,@      &@      &@      $@               @     �T@      n@      @      $@     @b@      2@     ��@     �D@     `{@      \@      @              5@     �T@                      9@      @      q@      "@      a@      7@       @              2@      T@                      8@      @      l@      "@     @[@      5@       @              *@     �B@                      (@             �f@      @     �J@      @       @              @     �E@                      (@      @     �F@      @      L@      ,@                      @       @                      �?             �H@              ;@       @                                                                      <@              &@       @                      @       @                      �?              5@              0@                       @     �N@     �c@      @      $@     @^@      &@     0t@      @@     �r@     @V@      �?              C@      `@      @      @     �N@       @     @q@      $@     �k@     �K@      �?              *@      Y@       @       @     �D@      @     �e@      @      d@      =@                      9@      <@      @       @      4@      @     @Y@      @     �O@      :@      �?       @      7@      >@      �?      @      N@      @     �G@      6@     �S@      A@               @      �?      @              @      &@      �?      @      @      (@      @                      6@      8@      �?             �H@       @     �D@      0@     �P@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJS�l-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?-!�FP<@�	           ��@       	                   �2@�cf���@+           0�@                           �?�t}�j@           �{@                          �1@��%��@L            �^@������������������������       �Z~�)�@.            �P@������������������������       ���쓎�@            �K@                           @�Zhc��?�            �s@������������������������       �\�a��s�?�            @n@������������������������       ����q@,             S@
                           �?N݄�@            ��@                          �7@ǁ8��@%            }@������������������������       �.�o!�P@�            �q@������������������������       ��ky��]@q             g@                           �?MU�u�@�             x@������������������������       �Rق��@v            `f@������������������������       �����p@�            �i@                           @�몹@�           z�@                           �?�q���4	@�           �@                           �?�[?^��	@�            �@������������������������       �\FZ�;@           �z@������������������������       �t��>H�	@�           ��@                           �?+mC�.@�            �w@������������������������       ����@             <@������������������������       �<���F@�            �u@                          �7@W�	�7@�           �@                          �3@n�Yu�4@           ��@������������������������       ��h�5�!@"           `|@������������������������       ���I
�@�            w@                          �<@��J�J�@�            �p@������������������������       �ʹ�5=W@�            �h@������������������������       �t5�DVR@*             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �s@     ȁ@      ;@      F@     P|@     �U@     ��@      l@     І@     �v@      :@             �Z@      h@      @      "@      Z@       @     �}@     �E@     �o@      V@      @              >@      H@              @      6@             `k@      @      U@      ;@                      *@      5@              @      $@              B@      @      ;@      "@                      @      0@                      $@              4@      �?      "@      @                      "@      @              @                      0@       @      2@       @                      1@      ;@                      (@             �f@      @     �L@      2@                      "@      6@                      @             �b@      �?     �E@      "@                       @      @                      @              @@      @      ,@      "@                     @S@      b@      @      @     �T@       @     p@      B@     @e@     �N@      @             �C@     �Q@      @      @      H@       @      c@      7@      T@     �A@      �?              1@      F@      �?      @     �B@      @     �Y@      (@      F@      ,@      �?              6@      ;@       @      @      &@      �?      I@      &@      B@      5@                      C@     @R@      �?              A@             @Z@      *@     �V@      :@      @              8@      B@                      7@              =@       @      A@      3@      @              ,@     �B@      �?              &@              S@      @      L@      @              4@     �i@     �w@      7@     �A@     �u@     �S@      �@     �f@     �}@     @q@      3@      3@      `@     �m@      1@      8@     `m@     �M@     �j@     �c@     �l@     `h@      1@      3@     �X@     `f@      1@      6@     �f@      G@     �`@     �\@     `d@     `d@      0@      @      3@      R@       @      &@      M@       @     @Q@     �C@     �R@      P@      @      .@      T@     �Z@      .@      &@     �^@      C@      P@     �R@      V@     �X@      (@              =@      M@               @      K@      *@     �T@      E@     �P@      @@      �?              @      @                      @      �?              $@      @       @                      :@     �J@               @     �I@      (@     �T@      @@      O@      >@      �?      �?     @S@     �a@      @      &@     �\@      4@     �v@      :@     �n@     @T@       @              F@     @^@      @      "@     �P@      1@     �r@      (@     �h@      H@       @              :@     �L@              @      ?@      @     �e@       @     �^@      ;@                      2@      P@      @      @      B@      ,@     �_@      @      S@      5@       @      �?     �@@      3@       @       @     �G@      @      P@      ,@     �H@     �@@              �?      8@      (@       @      �?      7@      @      K@      (@      G@      5@                      "@      @              �?      8@              $@       @      @      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�z�IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��W]@�	           ��@       	                     �?��ò��@�           �@                          �5@���`c@�           ��@                          �3@�'��@�             u@������������������������       ���NGZ@�            �h@������������������������       ��P�	3@W            `a@                           @O�ɄƮ	@�            v@������������������������       �華T�%	@�            @k@������������������������       �7O��E@T            �`@
                           @)�uֶ@�           `�@                            �?}����@^           ��@������������������������       �_o�:@�            �s@������������������������       ��N?�Z@�           ȃ@                           @ Vf�i+	@o            �@������������������������       �W/�Xp�@           P{@������������������������       ��e���[@P            �[@                          �4@Q��r�@<           ��@                           @+�]��n@N           0�@                          �1@��gL�@�            �m@������������������������       �ʼB�?/             T@������������������������       � Ӟ�<@^            �c@                           �?2����@�           ��@������������������������       �V M8X@�            w@������������������������       �Q�:�~�@�            pt@                            �?�� =)@�           ��@                          �5@����;@            �z@������������������������       ��|�3l�@9            �X@������������������������       �YWj^K�@�            `t@                           @�p?`�@�             w@������������������������       ����@�            �s@������������������������       �m��m~@              K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@     p�@      >@     �I@     0~@      V@     8�@      l@     Ј@     0v@      :@      4@     �g@     `u@      4@      B@     �t@     @P@     �w@     �g@     �u@     �n@      0@      @     �J@      \@      @      0@     �X@      2@     �`@      R@     �^@     �J@      @              .@     @P@               @      F@      "@     @S@      <@     �R@      7@                      @     �A@                      0@      @      K@      7@     �G@      ,@                      $@      >@               @      <@      @      7@      @      <@      "@              @      C@     �G@      @      ,@      K@      "@     �K@      F@     �G@      >@      @      @      6@      =@              @      =@      "@      G@      0@      A@      1@      @              0@      2@      @      @      9@              "@      <@      *@      *@      �?      .@     @a@     �l@      .@      4@      m@     �G@     @o@     �]@     @l@     @h@      &@      @     �U@     �`@      $@      (@     �a@      ;@     �h@      G@     `d@     �^@      @              :@      A@      @      @     �C@      (@     �M@      (@     �R@     �I@              @     �N@     �X@      @      @     �Y@      .@      a@      A@     @V@      R@      @      &@     �I@     @X@      @       @     �V@      4@      K@      R@     �O@     �Q@      @      @     �D@     @S@      @       @     �Q@      *@     �E@     �H@     �K@     �P@       @      @      $@      4@                      4@      @      &@      7@       @      @      @             �W@      o@      $@      .@      c@      7@     H�@      A@     �{@      [@      $@              K@     �^@      @      @     �M@      �?     �x@      *@     @l@     �H@      �?              8@     �H@                      .@      �?     @X@       @      C@      @                      @      $@                      �?              J@       @      &@      �?                      5@     �C@                      ,@      �?     �F@      @      ;@      @                      >@     �R@      @      @      F@             �r@      @     �g@     �E@      �?              $@      @@       @      @      =@             �f@      @     @T@      6@                      4@      E@      �?      �?      .@             �]@      �?     �Z@      5@      �?              D@     @_@      @       @     �W@      6@     `g@      5@     �k@     �M@      "@              9@     @S@      @      @      @@      3@      W@      .@      ^@     �B@      �?                      A@                       @       @      :@      �?      8@       @      �?              9@     �E@      @      @      8@      1@     �P@      ,@      X@     �A@                      .@      H@      @      @      O@      @     �W@      @      Y@      6@       @               @     �A@      @      @     �I@      @     @V@      @     �W@      5@                      @      *@      �?              &@              @       @      @      �?       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�HdhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?&��su@�	           ��@       	                    �?|���X	@�           ܘ@                          �5@��ǘ@)           �}@                           �?C]�<��@�             m@������������������������       �Y��y�@@            @Y@������������������������       �����@U            ``@                            �?��,���@�             n@������������������������       �V�I0��@-             R@������������������������       ���1���@g             e@
                           @)s����	@�           |�@                           �?W=N]^q	@�           ��@������������������������       �'��D0t@�            �q@������������������������       ��Xx��	@           �y@                          �:@���7�	@           0z@������������������������       �^/�m�	@�             t@������������������������       ����@=            @X@                           �?�-"��@�           $�@                           @�Uz� @�           H�@                          �;@"�I��@l            �d@������������������������       ��EpD�@`             b@������������������������       ���t@             4@                          �4@��8�O=@o            �@������������������������       �c8N��1�?�            �v@������������������������       �k��u�@�             k@                           @�3��@�           ��@                           �?N��s��@\           ��@������������������������       �����@?             [@������������������������       �AV(�@            �@                          �2@:�cd�@x            �g@������������������������       ���?
��?             =@������������������������       �w%	gc@g             d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     0s@     `�@      A@      O@     @|@      U@     ��@     �k@     ��@      w@      7@      9@      h@     @l@      7@      =@     �n@      F@     @i@      a@      o@     �h@      3@      �?      L@      Q@      �?      @     �O@      @     @X@     �@@     �X@     �E@      �?              .@      ?@      �?      @      5@      @     �Q@      0@     �I@      4@                       @      0@                      @             �D@      @      >@      @                      *@      .@      �?      @      0@      @      =@      (@      5@      1@              �?     �D@     �B@               @      E@      �?      ;@      1@      H@      7@      �?      �?      0@      $@                      .@      �?      $@       @      .@      �?      �?              9@      ;@               @      ;@              1@      .@     �@@      6@              8@      a@     �c@      6@      8@      g@     �C@     @Z@      Z@     �b@     �c@      2@      ,@     �T@     �X@      0@      "@      \@      9@      R@      E@     �\@     @Z@      $@       @      9@     �D@      @      @      I@       @      H@      1@     �I@      A@       @      (@      M@     �L@      $@      @      O@      1@      8@      9@     �O@     �Q@       @      $@     �J@      N@      @      .@      R@      ,@     �@@      O@     �A@     �I@       @      @     �E@     �J@      @      ,@     �L@       @      <@      H@      <@      8@      @      @      $@      @              �?      .@      @      @      ,@      @      ;@      �?             �\@     �t@      &@     �@@     �i@      D@     X�@      U@     0�@     `e@      @              8@     @W@      �?      @      G@      &@     �u@      &@     �e@      @@      �?              "@      $@              @      .@       @     �P@      @      E@      $@      �?               @      "@              @      $@       @     �P@      �?      B@      "@                      �?      �?                      @                      @      @      �?      �?              .@     �T@      �?      @      ?@      "@     `q@      @     �`@      6@                      &@      E@              @      3@              i@      @     �R@      $@                      @     �D@      �?              (@      "@     �S@       @     �L@      (@                     �V@     �m@      $@      :@     �c@      =@      }@     @R@     �u@     `a@      @             �P@     @j@       @      8@     �b@      9@     `z@     �J@     �s@      \@                      @      *@              &@      *@      @      .@      *@      1@      ,@                     �N@     �h@       @      *@      a@      3@     py@      D@     �r@     �X@                      8@      ;@       @       @      $@      @      F@      4@      :@      ;@      @                      @              �?                       @              @      (@                      8@      6@       @      �?      $@      @      B@      4@      7@      .@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�(?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�ŭ_@�	           ��@       	                    �?t%��C=@�           �@                           @�$���=@�           (�@                          �7@�4�4�p@�            `v@������������������������       ��K:)@�             o@������������������������       ����6�@I            �[@                          �5@[�l��}�?�            �o@������������������������       �_���I�?u            �e@������������������������       ��>=���@4            @T@
                           �?��ٯ�@j           ��@                          �<@��K��@�            `p@������������������������       ���0F��@�            �l@������������������������       �saW@             A@                            @p���� @�            �t@������������������������       �XJ4v@�            @q@������������������������       �g�1�1�?$             M@                           @���vT@�            �@                          �1@D�����	@�           ��@                            @a��uw@j            `f@������������������������       ��%R{m@A             \@������������������������       �����#�@)            �P@                           �??�����	@\           ��@������������������������       �.�J�6
@�           $�@������������������������       �$��;/@�            Pv@                            �?�Ö���@�           ��@                          �;@�"���@�            �p@������������������������       ��~��;@�            @n@������������������������       ���K����?             6@                          �7@�����@1           8�@������������������������       �V�d\�@�           �@������������������������       �`�.;	@�            @m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     ��@      D@      J@     P{@     @T@     �@      i@     �@     �u@      C@      �?      U@     �c@      @      &@      T@      *@     �|@      C@     �q@      S@      @      �?     �D@     @S@       @      $@     �A@      (@     pp@      5@     @\@      B@       @      �?      B@     �F@       @      @      :@      "@     �]@      0@     @P@      ?@       @              4@      ;@              �?      8@      "@     @X@      &@      E@      .@       @      �?      0@      2@       @      @       @              6@      @      7@      0@                      @      @@              @      "@      @      b@      @      H@      @                      @      .@              @      @             �\@      �?      <@      @                      �?      1@                      @      @      =@      @      4@       @                     �E@     �S@      �?      �?     �F@      �?     �h@      1@      e@      D@      @             �A@     �D@              �?     �@@              G@      $@     �Q@      7@       @              ?@     �B@                      :@             �F@       @     �P@      (@       @              @      @              �?      @              �?       @      @      &@                       @      C@      �?              (@      �?      c@      @     @X@      1@      �?              @     �B@      �?              "@      �?      \@      @     �U@      0@      �?              �?      �?                      @              D@      �?      &@      �?              6@      k@      z@     �B@     �D@     Pv@      Q@     ��@     `d@     @�@     �p@     �@@      5@     `d@      p@      >@     �@@      o@      J@     �h@      a@     �k@     �f@      =@      �?      4@      A@      @              &@      �?     �E@       @     �@@      7@              �?      @      9@                      @      �?      =@       @      3@      1@                      *@      "@      @              @              ,@              ,@      @              4@     �a@      l@      9@     �@@     �m@     �I@      c@      `@     �g@     �c@      =@      4@     �]@     �c@      7@      9@     `g@      B@     �X@     �Y@      `@      \@      ;@              8@      Q@       @       @      I@      .@     �K@      ;@     �N@     �F@       @      �?      K@     �c@      @       @     @[@      0@     �v@      :@     �r@     �V@      @              ,@      ?@                      8@      @     �W@      "@     �Q@      3@                      *@      :@                      8@      @     �W@      "@     �N@      (@                      �?      @                                                      "@      @              �?      D@     �_@      @       @     @U@      *@     �p@      1@     �l@     �Q@      @              6@      Z@      @      @      H@      "@     �k@      @      e@     �G@      @      �?      2@      7@      @      @     �B@      @     �H@      (@     �M@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJR�4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��v�f\@�	           ��@       	                   �;@�z��@�           ��@                           �?�$B�7@�           ��@                           �?���/�@v           ��@������������������������       �s�ڐ��@            |@������������������������       �~�|@cg@e            �c@                           @�s*�@U           �@������������������������       �����s@�           ��@������������������������       �v���(	@c            @d@
                           �?�&�u��	@�            �s@                            @�$��@R             a@������������������������       �xb���/@0            �S@������������������������       ���\�@"             M@                           �? &�`p�	@n            �f@������������������������       ��E��u@!             K@������������������������       �,����	@M            �_@                            �?�n�iO#@           ��@                          �5@=8�B��@�            `v@                          �1@��y���?�            �l@������������������������       ���R�?1            �R@������������������������       ���:���?`            @c@                           �?��~@T            @`@������������������������       ��G�*�@)            �M@������������������������       ��j��@+            �Q@                          �4@�rL@5           �@                          �1@w ����@�           ��@������������������������       �d)�x;.�?�             p@������������������������       ���	YjB@           {@                           @v:�dP@�           ��@������������������������       �(��X!Y@           �x@������������������������       �\N1��<@�            `i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     H�@     �A@      P@     �|@     �V@     `�@      m@     ��@     �r@      A@      &@     @l@     Pu@      6@     �G@     Pt@     �Q@     @x@     �g@     `y@      k@      :@      @      h@     �r@      4@     �@@     �q@     �F@      w@     �b@     `w@      c@      8@             �M@     @U@      @      &@     @Q@       @     �c@      =@     �b@      @@      @             �F@     �Q@      @      $@      K@      �?      Y@      <@     �Y@      ;@      @              ,@      ,@              �?      .@      �?      M@      �?     �G@      @              @     �`@     �j@      ,@      6@      k@     �E@     �j@     �^@      l@     @^@      5@       @      ^@     �g@      *@      5@      h@      B@     �h@      V@     �j@     @Z@      *@      @      *@      ;@      �?      �?      9@      @      .@      A@      (@      0@       @      @      A@     �D@       @      ,@     �C@      9@      2@      D@      @@     �O@       @      @      $@      7@      �?      @      7@      &@       @      *@      2@      =@                      @      "@      �?              "@      "@       @      $@      (@      3@              @      @      ,@              @      ,@       @              @      @      $@              @      8@      2@      �?      &@      0@      ,@      0@      ;@      ,@      A@       @       @      @      @                       @      @      @      @      @      $@              �?      2@      (@      �?      &@       @       @      "@      5@      &@      8@       @       @      S@     �j@      *@      1@     �`@      5@     @�@      E@     `z@     @T@       @              .@      A@      @              6@      @     �d@      .@     �R@      3@                      @      3@                      *@             �`@      @      H@      @                              @                      @             �H@              "@      @                      @      *@                       @             @U@      @     �C@      �?                      $@      .@      @              "@      @      @@      (@      ;@      *@                      @      @                      @      �?      0@      @      (@      @                      @       @      @              @      @      0@      @      .@      @               @     �N@     @f@       @      1@      \@      ,@      |@      ;@     �u@      O@       @              B@      Z@      @      $@      @@      @     �q@      *@      f@      ;@      �?              @     �C@              @       @              _@      �?     �Q@      @      �?              ?@     @P@      @      @      8@      @     �c@      (@     �Z@      7@               @      9@     �R@       @      @      T@      &@     @e@      ,@     @e@     �A@      @       @      0@      G@              @     �J@      @     �`@      @     @Z@      0@      @              "@      <@       @      @      ;@      @      B@       @     @P@      3@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJi�EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��%�D@�	           ��@       	                    �?K�6���@\           �@                           �?H��=@�           @�@                            �?%�<�[~@	           �z@������������������������       �+�LN�@:            �V@������������������������       �)�i� �@�            0u@                           @IP�}�@�            �u@������������������������       �b�xS��@|            �f@������������������������       ����� @b            �d@
                          �1@ ��&�@u           ��@                           �?�t�Pl@�            w@������������������������       ����@A            @X@������������������������       ��J��CK@�             q@                           �?ܤ�m@�           4�@������������������������       ���4 �j@5            �U@������������������������       �9n�Y�`@T           ��@                           �?��7��@B           �@                           �?���=Dc@�           ��@                            �?פ�&��	@�            �r@������������������������       ��_(1v@c            �a@������������������������       ����G
@f            �c@                           @��r��5@
           �|@������������������������       �O8P�E@@            @]@������������������������       ��Hxk}@�            @u@                           �?p^�2�@o           `�@                          �7@�z��	@T           ��@������������������������       �5ѐe��@X             b@������������������������       �x��܇�	@�            Px@                          �>@Z����@           p{@������������������������       �)#p�r@           Py@������������������������       ���A6�@             A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     X�@      A@     �O@     0{@      U@     Ў@     �g@     P�@     Pv@      >@      @     @^@     �u@      $@      =@     �h@      >@      �@     �U@      �@      c@      (@              F@     �^@      �?      @     �E@      @     �r@      4@     �g@     �E@      �?              3@     �Q@      �?      @      <@      @     �e@      *@     �V@      6@      �?                      3@               @      @       @      D@      @      2@      @                      3@      J@      �?      @      8@       @     �`@      $@     @R@      3@      �?              9@      J@               @      .@             �_@      @     @X@      5@                      0@      7@               @      &@              H@      @     �M@      3@                      "@      =@                      @             �S@      @      C@       @              @     @S@      l@      "@      6@     �c@      :@      w@     �P@     �t@     �[@      &@      �?      3@      K@      �?       @      <@              a@      &@     @W@      7@              �?      @      2@      �?      �?      .@              *@      @      9@      .@                      ,@      B@              �?      *@              _@       @      Q@       @              @      M@     `e@       @      4@      `@      :@      m@      L@     `m@     �U@      &@      @       @      .@              �?      (@       @      @      @      @@      "@              �?      L@     �c@       @      3@      ]@      8@     `l@      J@     `i@     �S@      &@      *@     �d@     �m@      8@      A@     �m@      K@     �s@      Z@     `t@     �i@      2@      @      O@     �Z@      (@      3@     �Y@      0@      c@     �B@     �a@     �X@       @      @      :@     �J@      $@      &@      E@      $@     �A@      5@      >@     �J@      @      �?      (@      6@      @      @      4@              3@      0@      $@      @@      @      @      ,@      ?@      @      @      6@      $@      0@      @      4@      5@      @              B@      K@       @       @     �N@      @     @]@      0@     �[@     �F@      �?              *@      $@               @      5@      @      9@      "@      8@      "@      �?              7@      F@       @      @      D@      @      W@      @     �U@      B@              "@     �Y@     �`@      (@      .@     �`@      C@     @d@     �P@      g@     �Z@      $@      "@     @P@      T@      &@      "@     �S@      0@      O@      F@     �T@     @P@      $@      @      @@      9@      @      @      0@       @      @      "@      >@      ,@              @     �@@     �K@      @      @     �O@      ,@     �L@     �A@     �J@     �I@      $@              C@      J@      �?      @      K@      6@      Y@      7@     �Y@     �D@                      C@      J@      �?      @     �D@      6@     @W@      4@     �W@      C@                                              �?      *@              @      @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJn֙yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��Z�"@@�	           ��@       	                    �?�*<NT�@X           �@                           �?�"�7+	@�           �@                           �?N�	T@&           �|@������������������������       �ִwG�x@�            �h@������������������������       ���E�@�            �p@                          �:@,�m7/�	@�           ��@������������������������       ��@�D�W	@4           ؋@������������������������       �\�!�j�	@�             n@
                          �1@��
	Ft@`           ��@                          �0@�.� @:            �X@������������������������       ��-�l@            �A@������������������������       �F��* @&             P@                            �?n��^�@&           0}@������������������������       �$���>@�            �p@������������������������       ���E@z             i@                           @ǯCI��@?           d�@                           �?=:T���@�           ��@                           @o����?�            �y@������������������������       �7O�"� @�            �p@������������������������       �;	/��8�?V            @b@                           �?���
�E@�           `�@������������������������       ��AhM��@            �E@������������������������       ��U�c�@�           �@                            @��8yHv@U           ��@                          �;@	�f�@�             z@������������������������       ��`Њ�@�            �v@������������������������       ��I�,$@            �L@                           @�4� @V            �a@������������������������       ��$W�i @+            @Q@������������������������       �����@+            @R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �s@     Ȁ@      8@      F@     `|@     �U@      �@     �j@     ��@     �u@      @@      9@     �k@      t@      5@     �@@     �s@      O@     �w@     `e@     �u@     `n@      :@      9@      e@     @o@      2@      6@      n@      G@     �l@     �^@     �o@     @h@      9@             �G@     �U@       @      @     �J@       @      [@      8@     �V@      F@       @              *@     �B@       @       @      3@       @     �K@      0@      <@      7@                      A@     �H@              �?      A@             �J@       @     �O@      5@       @      9@     @^@     �d@      0@      3@     �g@      F@     �^@     �X@      d@     �b@      7@      $@     �V@      b@      &@      1@     �b@      ;@      Z@     @R@     �a@     �Y@      4@      .@      >@      4@      @       @      C@      1@      2@      :@      4@     �G@      @              J@     �Q@      @      &@     �R@      0@     @b@      H@     �W@     �H@      �?              @      *@                      $@              H@      @      *@      @                       @      @                      @              *@              @      @                      �?      @                      @             �A@      @      $@       @                     �H@     �L@      @      &@     @P@      0@     �X@     �D@     �T@      F@      �?              ;@      ?@       @       @      B@      .@     �L@      3@      J@      3@      �?              6@      :@      �?      @      =@      �?     �D@      6@      >@      9@              �?     �W@      k@      @      &@     @a@      8@     ��@     �E@     0|@      [@      @      �?     �N@     ``@              @     �S@      0@     �~@      6@     �s@     @Q@      @              0@     �E@                      &@      @      l@       @      X@      .@                      *@      >@                      $@      @     �`@       @     �M@      ,@                      @      *@                      �?             �V@             �B@      �?              �?     �F@      V@              @     �P@      &@     �p@      4@      k@      K@      @      �?      @      "@              �?      @       @       @      @       @                             �C@     �S@              @      P@      "@     @p@      .@      j@      K@      @              A@     �U@      @      @      N@       @     `d@      5@     `a@     �C@      �?              ;@     �R@      �?      @     �I@       @      [@      .@     @Z@      8@      �?              6@      M@      �?      @      B@      @     �Z@      .@     @X@      0@      �?              @      0@                      .@      @       @               @       @                      @      (@       @       @      "@             �K@      @      A@      .@                      @      �?              �?       @             �B@      @      ,@      @                      @      &@       @      �?      @              2@              4@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @~���O@�	           ��@       	                   �2@�R\�&�@P           Ġ@                           �?��C�ԯ@/           �}@                           �?�5P�]�@g            �b@������������������������       ����/O!@*            �M@������������������������       �y��@=            @V@                           �?��
/�@�            Pt@������������������������       ���ɭE@N            �_@������������������������       ��}f5A @z            �h@
                          �8@�u$�Zs	@!           $�@                           �?/C�@�           �@������������������������       �f�d�8�@�            `r@������������������������       ���q	@�            �@                           �?0�M;\�	@�           �@������������������������       ����T,_@]             c@������������������������       ��c��+�	@,           �~@                           �?�7�.1@h           ��@                          �4@�A�w@�           ȃ@                            �?��S�8a�?�            @x@������������������������       �����?�            �j@������������������������       ��w%o�?r            �e@                            �?0O���D@�            �n@������������������������       �r��ZHc @"             J@������������������������       �B� �"b@|             h@                           @sLé]@�           ��@                           @�(�Z@�           4�@������������������������       ��Ė��@�           `�@������������������������       ���qf@�            t@                            �?*D�u�g@            �@@������������������������       ���1�@             1@������������������������       �+�%W�@	             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      s@     ��@      >@     �K@      }@     �U@     ��@     �l@     �@      u@      @@      ,@     �j@     �s@      9@      D@     pr@     �P@     Pw@     �g@     Pw@     �j@      <@             �C@     @R@              @     �L@       @     �a@      @@      U@      C@      �?              @      3@                      7@      �?     �K@      @      4@      .@      �?              �?       @                      @      �?      ?@      �?      @      @                      @      &@                      1@              8@      @      *@      &@      �?              @@      K@              @      A@      �?      V@      9@      P@      7@                      &@      .@              @      $@              G@      @      <@      "@                      5@     �C@                      8@      �?      E@      6@      B@      ,@              ,@     �e@     @n@      9@      B@     �m@      P@     �l@     �c@     r@      f@      ;@      @      [@     �c@      2@      :@      c@      8@     �c@     �P@     �i@     �W@      .@              2@      I@      �?       @     �C@      @      N@      .@     �K@      C@      @      @     �V@     �Z@      1@      2@     �\@      2@     @X@     �I@     �b@     �L@      &@      @     �P@     @U@      @      $@     @U@      D@     @R@     �V@     @U@     �T@      (@      �?      &@      1@      �?       @      4@      @      <@      *@     �@@      3@      @      @      L@      Q@      @       @     @P@     �B@     �F@     @S@      J@     �O@       @       @      W@     �k@      @      .@      e@      4@     H�@     �D@     �z@     @^@      @              5@     @S@              �?      D@      @     Pr@      $@     �c@      <@      �?              ,@      A@              �?      2@             @j@      @     �V@      .@      �?              @      4@                      ,@             �[@             �I@      (@                       @      ,@              �?      @             �X@      @     �C@      @      �?              @     �E@                      6@      @     �T@      @     �P@      *@                              @                      "@       @      :@              @       @                      @     �B@                      *@      @     �L@      @     �M@      &@               @     �Q@     �a@      @      ,@      `@      ,@     @v@      ?@     q@     @W@      @       @     �O@     �a@      @      (@     �^@      &@     v@      <@     �p@     �V@      @       @      G@     @Z@              @     �T@       @     0q@      .@     �g@     �L@       @              1@     �B@      @       @      D@      "@     �S@      *@     �S@      A@      �?               @      �?               @      @      @      @      @      @       @                      @                       @       @      @               @      @      �?                      @      �?                      @              @      �?      �?      �?        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ6�yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�F�)X@�	           ��@       	                    �?�M<��@Q           ��@                          �1@{��PDo@�           0�@                           �?�ܔ_Z� @�            Pp@������������������������       ���
�@P             _@������������������������       ������?Q             a@                           �?)Z�Q��@2           |@������������������������       ��+��>�@�             p@������������������������       ��b�"@�             h@
                           �?3D���@~           ,�@                           �?�wN�^=	@A           h�@������������������������       �?�<�32@�            �m@������������������������       ��>g�	@�            r@                          �4@��k:�@=           ��@������������������������       ���m*��@�           �@������������������������       �3r�"�@e             d@                           �?���P�@H           ��@                          �=@�f���@(           @                           �?��R��@�            0{@������������������������       �_�vi1x@z             i@������������������������       �X��Q��@�            @m@                          �?@#�p�z�@)             O@������������������������       ���H�@             @@������������������������       ��֬<��@             >@                           @,E�^�0	@            �@                           @��s��	@�           ��@������������������������       �� `:�	@�           0�@������������������������       ��
l*��@           �y@                            �?����4@j            �d@������������������������       �y�<P		@             �F@������������������������       �̥�c?@J            �^@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �q@     ��@      <@     @P@      |@     @U@     0�@     `n@     Љ@     `v@     �@@      @      \@     s@      $@      2@      k@      ?@     ��@      ]@      ~@      c@      &@             �A@     �S@                     �L@      @     �s@      8@     �d@      =@       @               @      9@                      7@             �a@      $@     �C@      *@      �?              @      *@                      ,@             �P@      @      $@      $@                      @      (@                      "@             �R@      @      =@      @      �?              ;@     �J@                      A@      @     @e@      ,@      `@      0@      �?              &@      9@                      7@      @      [@      (@     �O@      @      �?              0@      <@                      &@              O@       @     @P@      "@              @     @S@     `l@      $@      2@      d@      9@     @v@      W@     �s@     �^@      "@      @      C@      U@      "@      "@     �T@      ,@     @P@      K@     �V@      O@      "@              (@     �G@              @     �B@      @      B@      =@     �G@      0@      �?      @      :@     �B@      "@      @      G@      "@      =@      9@      F@      G@       @             �C@     �a@      �?      "@     @S@      &@     0r@      C@      l@     �N@                      B@      ]@      �?       @      P@      @     �n@     �A@     �e@      J@                      @      ;@              �?      *@      @      G@      @      J@      "@              @     @e@     �l@      2@     �G@      m@      K@     �t@     �_@     �u@     �i@      6@              E@      N@      @      "@      J@      @     @a@      <@     �[@      G@       @              C@     �L@      @      @     �C@      @      `@      2@     �Y@     �B@      �?              ?@     �A@       @      @      :@      �?      >@      ,@      D@      1@      �?              @      6@      @              *@      @     �X@      @      O@      4@                      @      @              @      *@              "@      $@       @      "@      �?                       @              @      @              @      @       @      @      �?              @      �?               @      "@               @      @      @      @              @      `@      e@      *@      C@     �f@     �H@      h@     �X@     @m@      d@      4@      @     �[@     @b@      "@      C@     �c@     �F@     `d@      R@      j@     @c@      ,@      @     �T@      V@      @      ;@      Z@     �C@     @R@      N@      \@     @Y@      ,@       @      ;@      M@      @      &@      J@      @     �V@      (@      X@     �J@                      2@      6@      @              9@      @      =@      ;@      :@      @      @              @      @      @              @      �?      @       @      "@      @      @              (@      3@      �?              5@      @      9@      3@      1@       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�M�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�	�0�.@�	           ��@       	                   �;@JF�?��@�           ��@                           �?,]�(Q?@�           `�@                           �?
L�Q{�@�           �@������������������������       �ҝMn�@�            r@������������������������       ��\�Zd	@<           �@                          �7@.���@�           ؑ@������������������������       ������@/           ��@������������������������       �
�{��@�            �q@
                           �?�V�aY�@�             s@                           �?�S���@1            �S@������������������������       �"[&��|@             :@������������������������       �J����@            �J@                           @��t		@�             l@������������������������       �Vɲ�P@D            @Z@������������������������       ����8	@P             ^@                           @h=H�@?           �@                          �7@��'�f�@�           0�@                            @_���~�@j           ��@������������������������       ��޶@$           @�@������������������������       ��D��BF�?F            @[@                           �?��/W�q@�            �j@������������������������       ��D�Z���?             F@������������������������       ���BH��@o            `e@                           �?���B@J           P@                            @�r;�ŧ@y            �f@������������������������       �aZ��@Z            @a@������������������������       �|�2,���?            �E@                          �;@�c�fԇ@�             t@������������������������       ���7^�@�            q@������������������������       �ϼ�M�@            �G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     8�@     �@@      N@     �{@     �S@     ,�@     `m@     �@     Pv@      4@      .@      i@     0u@      :@     �B@     t@      N@      y@     �h@     y@      m@      1@      *@     `d@      s@      5@      >@     pq@     �F@     �w@     �d@     pv@     �d@      0@      @      N@     `a@      0@      .@      \@      6@     `f@      P@     @\@     @Q@      "@              5@      F@      @      @      >@      @      Z@      3@      G@      *@              @     �C@     �W@      (@      &@     �T@      2@     �R@     �F@     �P@      L@      "@      "@     �Y@     �d@      @      .@     �d@      7@     �i@      Y@     �n@      X@      @      @     @U@      `@      �?      ,@      ]@      "@     `b@     �Q@     �h@     �T@      @      @      2@     �C@      @      �?     �I@      ,@     �L@      >@     �H@      ,@       @       @     �B@     �@@      @      @      E@      .@      3@      A@      E@     �P@      �?               @      @      �?      �?      @      �?      @      $@      4@      5@                      @      �?              �?      @              �?      @      @      @                      @       @      �?              @      �?      @      @      .@      0@               @      =@      >@      @      @     �A@      ,@      (@      8@      6@      G@      �?      �?      (@      $@       @       @      .@              @      0@      *@      ;@              �?      1@      4@       @      @      4@      ,@      @       @      "@      3@      �?      �?      T@     �j@      @      7@     @_@      3@     ȃ@     �B@      y@     @_@      @      �?      J@     �a@      �?      @     @R@      (@     �~@      2@     �q@     �T@      @             �A@     �^@      �?       @     �F@       @     �z@      @     `m@     �P@      �?             �@@     @\@      �?       @      D@      @     �w@      @     �g@     �P@                       @      "@                      @       @     �F@              F@      �?      �?      �?      1@      5@              @      <@      @     �O@      &@     �H@      .@       @              �?      @                              @      5@              $@      �?              �?      0@      ,@              @      <@              E@      &@     �C@      ,@       @              <@     @Q@      @      1@      J@      @      b@      3@      ]@     �E@                       @      >@      �?      �?      ,@             �Q@      @     �F@      @                      @      =@      �?              ,@              H@      @     �@@      @                       @      �?              �?                      7@       @      (@       @                      4@     �C@      @      0@      C@      @     @R@      ,@     �Q@     �B@                      .@      @@      @      *@      ?@      @     �Q@       @     �P@      ;@                      @      @       @      @      @      �?       @      @      @      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�D�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�K��3@�	           ��@       	                    �?@ugA=�@�           p�@                           �?h�7��@"           �|@                           �?D��L�E@S             a@������������������������       �8sO�d@"            �L@������������������������       ���Fý@1             T@                           �?����9	@�            t@������������������������       ����U��@D             [@������������������������       ����4`	@�            �j@
                           �?7����@u           ��@                           @���}�@�            r@������������������������       ��� �@s            `f@������������������������       �J��O�K@?            �[@                          �5@+��@�            s@������������������������       �Lr�h��?y             g@������������������������       ����@J            @^@                           �?�X�ֲA@'           Z�@                           �?�'&LI	@�           �@                          �3@���w5	@            �|@������������������������       �(�P�N'@P            ``@������������������������       ��O1��	@�            �t@                           @�p�tu	@�           ȅ@������������������������       ��9`�+�@S           ��@������������������������       ��a6N�@j             e@                           @Dc��1�@J           ��@                            @�P�s�\@�           P�@������������������������       ��FVb=�@2            }@������������������������       �?���@�            @k@                           �?#i,�Ah@�           ��@������������������������       ��(�9�� @�            Pv@������������������������       �����C@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     p�@      :@     �M@     �z@     �P@     �@     `j@     ��@      t@      E@      @     @S@     �b@      @      &@      ^@      9@     `t@     �L@     @g@     �R@      2@      @     �F@     �Q@      @       @     �R@      (@      T@     �D@     �R@      ;@      1@       @      1@      2@                      .@      @      @@      @     �@@      (@               @      @      $@                      $@              3@      �?      "@      @                      ,@       @                      @      @      *@      @      8@      "@               @      <@     �J@      @       @      N@      "@      H@      B@      E@      .@      1@              @      ?@      @              6@       @      *@      *@      $@      @      @       @      7@      6@               @      C@      @     �A@      7@      @@      &@      (@              @@     �S@      �?      @     �F@      *@     �n@      0@     �[@      H@      �?              "@      D@              �?      ;@       @     �]@      @      O@      8@                      @      ?@              �?      &@             �R@      @     �A@      1@                      @      "@                      0@       @      F@              ;@      @                      7@      C@      �?       @      2@      &@      `@      $@     �H@      8@      �?              @      9@                      @      @     @Z@       @      @@      @                      4@      *@      �?       @      &@       @      7@       @      1@      1@      �?      3@      l@     �{@      6@      H@     `s@     �D@     ��@     @c@     ��@     �n@      8@      2@     �^@     �h@      (@      ;@      e@      ;@      d@      V@     `f@     @a@      5@      @      H@      T@      "@      &@     �R@      ,@     @Q@      7@     �L@     @P@      @       @      @      1@                      9@      @      C@       @      0@      0@              @     �E@     �O@      "@      &@     �H@      $@      ?@      .@     �D@     �H@      @      (@     �R@     @]@      @      0@     �W@      *@     �V@     @P@     �^@     @R@      .@      @     �P@      S@       @      *@     @Q@      *@     �S@     �E@     �Y@      L@      @      @      "@     �D@      �?      @      :@              (@      6@      3@      1@      &@      �?     �Y@     �n@      $@      5@     �a@      ,@     ��@     �P@     P|@     �Z@      @      �?     @P@     @Y@      �?      @     �S@      &@     �e@     �A@     `c@      I@      @      �?     �F@      Q@      �?      @     �M@      &@     @X@      7@     �]@     �@@       @              4@     �@@              �?      4@             �S@      (@      B@      1@      �?             �B@     �a@      "@      .@      O@      @     �v@      ?@     �r@     �L@                      "@      M@               @      *@              c@      0@     �X@      @                      <@     @U@      "@      *@     �H@      @     �j@      .@     �h@      I@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ϳ'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����X@�	           ��@       	                    �?,U@���@           ��@                          �6@Ns�c0@�           @�@                          �0@M�@           �|@������������������������       ��8' @$            �R@������������������������       ��ΰ��@�            @x@                            @�lH���@v            @g@������������������������       ��p�y^@N            �_@������������������������       ��@�@(            �M@
                          �5@���s�@�           ��@                          �2@��<m3V@�            w@������������������������       �[�ʓ�@}            �h@������������������������       ���7�B�@m            �e@                          �>@&��鬋@�            `m@������������������������       �s�4D�E@�            �j@������������������������       ������ @             5@                           @dH��4@�           ʤ@                           @�[r�@�           �@                          �2@>�#	@`           �@������������������������       �7����@�             r@������������������������       �����]�	@�           ��@                          �7@���.A�@\           X�@������������������������       ��a�@�           ��@������������������������       ��˜��@�            `n@                           �?E�ů	@�            `u@                           �?pVhP��@C            �Y@������������������������       ��n,��@             K@������������������������       � �9?�.@$            �H@                          �<@]�x	@�            �m@������������������������       �Bd�@~            �h@������������������������       ���@            �D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@      t@     ��@      8@     �P@      |@      R@     ��@      n@     �@      u@      ?@      �?     �V@     `f@      @      .@     �Z@      .@     �|@     �@@      q@      Q@      @      �?     �D@     �T@      @      (@      J@      $@     �q@      6@     �Y@      B@                      4@      K@              "@      B@      @      n@      (@     @P@      4@                              @                      .@              C@      @      @      @                      4@     �G@              "@      5@      @     @i@      "@      M@      0@              �?      5@      =@      @      @      0@      @      F@      $@      C@      0@              �?      2@      8@                      @      @      8@      @      =@      ,@                      @      @      @      @      $@              4@      @      "@       @                      I@      X@      �?      @      K@      @      f@      &@      e@      @@      @              8@      M@              @      6@              a@       @     �Z@      .@       @              $@      4@              @      *@             �V@       @      H@       @       @              ,@      C@                      "@             �G@              M@      @                      :@      C@      �?              @@      @      D@      "@     �O@      1@      @              8@     �A@      �?              7@      @      B@      @     �O@      1@      @               @      @                      "@              @      @                              4@     �l@      v@      3@      J@     �u@     �L@     ��@      j@     h�@     �p@      9@      *@     �g@     �s@      0@     �G@     �r@     �E@     P@     �c@     @~@     `m@      0@      (@      b@     @g@      .@      A@     �h@      @@     @h@     ``@     `l@     �c@      0@      @      .@      D@              �?      E@             �R@     �@@      H@      ?@              "@     @`@     @b@      .@     �@@     `c@      @@     �]@     �X@     `f@      `@      0@      �?      F@     �`@      �?      *@     @Y@      &@     0s@      <@     p@      S@                      ?@     @\@      �?      @     �K@      &@     Pp@      *@     �g@      H@              �?      *@      3@              @      G@              G@      .@      Q@      <@              @      D@      A@      @      @      G@      ,@     �N@     �H@     �D@     �@@      "@              3@      $@       @       @      0@      $@      *@      3@      @      @       @              &@      @       @              $@       @              &@      �?      @      �?               @      @               @      @       @      *@       @       @      �?      �?      @      5@      8@      �?      @      >@      @      H@      >@      C@      :@      @      @      0@      7@      �?      @      4@      @      H@      6@     �A@      1@      @      @      @      �?                      $@      �?               @      @      "@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ&�|hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����|Z@�	           ��@       	                    �?�ҕ!�@           ؓ@                           �?֋��$�@�           ��@                           �?e�b�X@�            �j@������������������������       ��D=�3@=            @T@������������������������       � `���@S            �`@                           @���!\@            z@������������������������       �ܽ�w@k            �d@������������������������       ��2�ŷ @�            `o@
                          �<@\3�`�@�           �@                          �1@�$!@f           X�@������������������������       ��F�1Q��?R            �`@������������������������       �����@           p|@                            @FR(fdY@             K@������������������������       �+z����@             E@������������������������       ��D=�U��?             (@                           @�z��E@�           ��@                           �?Qr��v	@�            �@                           @��H�	@�           �@������������������������       �VaX��	@�           ��@������������������������       ����Lj�@             ;@                          �2@��bֿ@           Px@������������������������       ��N�6�@@             W@������������������������       �iɞ̝o@�            �r@                            �?�E�P�=@�           ,�@                           @���~��@�            @n@������������������������       �7rOy��@S             `@������������������������       ������@N            �\@                           @�����|@7           Ȍ@������������������������       ��JŲÊ@�           �@������������������������       ���1��@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �q@     8�@      6@      M@     @}@     �X@     ��@     `j@     �@      w@      <@      �?     �Q@     �e@      �?      *@     �\@      1@     `z@      H@     `t@     �T@       @      �?      <@      S@      �?      (@     �J@      .@     �m@      =@     @a@     �B@       @      �?      0@      9@      �?      &@      6@      @      I@      7@     �C@      3@       @      �?       @      @                      ,@              5@      @      4@      @                       @      2@      �?      &@       @      @      =@      2@      3@      ,@       @              (@     �I@              �?      ?@      &@     `g@      @     �X@      2@                      @      2@                      .@      &@     �P@       @     �C@      @                      @     �@@              �?      0@              ^@      @      N@      (@                      E@     �X@              �?     �N@       @      g@      3@     �g@     �F@                      D@     @V@                      H@       @     �f@      (@     �f@      @@                      �?      2@                       @              O@      �?      B@      @                     �C@     �Q@                      D@       @      ^@      &@     @b@      :@                       @      "@              �?      *@              @      @      @      *@                      �?      "@              �?      @              @      @      @      $@                      �?                              @                       @              @              2@     �j@     �y@      5@     �F@      v@     �T@     `�@     `d@     p}@     �q@      :@      0@     `a@      m@      (@     �A@     �n@     �P@     �g@     @`@     `h@      h@      9@      0@     @\@     �d@      &@      ;@     �h@      K@     �[@     �W@     �`@     �b@      8@      *@      \@     @d@      &@      ;@     �g@      K@     �[@      W@     �`@      b@      0@      @      �?       @                      @                      @      �?      @       @              :@     @Q@      �?       @     �I@      *@     �S@     �A@      O@      F@      �?              �?      5@                      @             �A@       @      0@      @                      9@      H@      �?       @      G@      *@      F@      ;@      G@      C@      �?       @     @R@      f@      "@      $@     �Z@      .@     �v@     �@@     @q@     �W@      �?              0@      @@      �?              .@       @     �X@      @      F@      ;@                      "@      5@      �?               @             �L@      @      ,@      .@                      @      &@                      @       @     �D@      @      >@      (@               @     �L@      b@       @      $@      W@      *@     �p@      :@      m@     �P@      �?       @     �C@     �[@       @      @     �L@      @     �i@      .@     �c@      C@      �?              2@      A@      @      @     �A@       @      P@      &@     �R@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�{83hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?F4�*�)@�	           ��@       	                     �?�
H��/@           x�@                          �8@�D��P�@�            �t@                           �?j�f�0|@�            �o@������������������������       ����T7@L            �_@������������������������       �t1��� @S             `@                          �<@٫�%��@*            �R@������������������������       �ÿ�7�@"            �N@������������������������       �V@���@             *@
                          �<@��CzS@E           ��@                           �?�H��@           ��@������������������������       ��I��Dd@�            pr@������������������������       ��.�G?\@a           h�@                            �?������@,            �P@������������������������       ����T��@             ;@������������������������       ����@            �C@                          �5@Õ��"@�           ֤@                           @�FX\�@}           �@                          �1@�p��j@>           ��@������������������������       �
���.�@�            �l@������������������������       �5�,@�           ��@                           @?��
@?           h�@������������������������       �6��Ɍ�@-            @������������������������       ��pՁ@             =@                           �?�rB� 	@           ��@                           @bM����	@�           ��@������������������������       ��[�4)
@�            Pw@������������������������       ��bf�N�@�            �l@                           @W��k�R@�           X�@������������������������       ��fp,�@7           �~@������������������������       �Rd��Д@[            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     (�@     �B@      H@     �}@     @T@     �@     �l@     ��@      t@      ;@              S@     �f@       @      "@     @[@      "@     p}@      H@     �p@     �Q@      @              ,@     �I@               @      >@      @     @_@      &@      S@      ,@       @              @      B@               @      8@      �?     �\@       @     �M@       @      �?              @      ,@               @      1@      �?      P@      @      4@      �?                      @      6@                      @             �I@      @     �C@      �?      �?               @      .@                      @       @      $@      @      1@      (@      �?               @      "@                      @       @      $@       @      .@      &@                              @                       @                      �?       @      �?      �?              O@     @`@       @      @     �S@      @     �u@     �B@     �g@      L@       @             �J@     �^@       @      @      R@      @     u@      <@     `g@     �C@       @              =@     �J@       @       @     �D@      @     @R@      0@      L@      3@      �?              8@     �Q@              �?      ?@      @     �p@      (@     ``@      4@      �?              "@      @              @      @              "@      "@      @      1@                      @      �?               @      �?              @      @       @      $@                      @      @               @      @              @      @       @      @              ,@     �i@      y@     �A@     �C@     �v@      R@     p�@     �f@     P�@     �o@      7@      @      S@      l@      &@      9@      e@      7@     pw@     �R@     �s@     @Y@      *@      @     �I@     @a@       @      2@      _@      $@     `l@     �C@     �i@     �N@      �?              @      C@       @      �?      7@             �T@      $@      L@      &@              @      F@      Y@      @      1@     @Y@      $@      b@      =@     �b@      I@      �?       @      9@     �U@      @      @      F@      *@     �b@     �A@     �[@      D@      (@              7@     @U@      @      @      F@      &@     �a@     �A@     �Y@      A@      &@       @       @      �?              �?               @      @              @      @      �?       @     ``@      f@      8@      ,@     �h@     �H@     �f@     �Z@     �i@     �b@      $@      @      R@      W@      1@      &@     �W@     �@@      P@     �P@     �M@     @T@      $@      @      K@      I@      ,@      "@     �L@      ;@      C@      ;@      A@      K@      @      �?      2@      E@      @       @     �B@      @      :@     �C@      9@      ;@      @      @     �M@      U@      @      @     �Y@      0@     �]@      D@     `b@     �Q@              @     �F@     �P@              @     �T@      "@     �Z@      >@     �Z@     �E@                      ,@      2@      @              4@      @      *@      $@      D@      ;@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�h��e'@�	           ��@       	                    �?P�� 	@�            �@                            @|����@*           �}@                           �?���f�@�            @q@������������������������       ����RS@P            �^@������������������������       �=�@a            @c@                           �?�9LF�@y            �h@������������������������       �C�2(@8            �W@������������������������       ����T0@A            @Y@
                           �?�=%��	@�           ��@                           �?>0���@=             Z@������������������������       �8�2@@             9@������������������������       �j����@-            �S@                           �?�t#��	@�            �@������������������������       ��� }Y*@�            �w@������������������������       �9+/�	@�           �@                           �?X�]I��@�           �@                           �?��5V6@�           ��@                            �?+��(>@            �x@������������������������       ���ο��@�            �k@������������������������       ��_��m�?o            �e@                          �8@Mv�g @�            Pu@������������������������       �u���Z��?�            �r@������������������������       ���B/@             �F@                           @���@�           ��@                           �? �.I�@           Pz@������������������������       ����E�@             A@������������������������       �dK�u ]@�            0x@                           @9�Վ�>@�           �@������������������������       ���l�@�           ��@������������������������       �>�0@             B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@      �@      >@      J@     `|@     �S@     �@     �j@     ؈@     �u@      ;@      ,@      f@      o@      6@      =@     �m@      G@     �m@      `@     �n@     `h@      5@             �M@      T@       @      @     @P@       @     �Y@      9@      T@      G@      @             �@@      E@       @       @     �C@       @      J@      4@      H@     �@@      @              (@      4@       @       @      4@       @      7@      $@      $@      4@      �?              5@      6@                      3@              =@      $@      C@      *@       @              :@      C@              @      :@             �I@      @      @@      *@                      $@      &@              @      .@              >@      @      2@      @                      0@      ;@              �?      &@              5@       @      ,@      "@              ,@     @]@      e@      4@      6@     �e@      F@     �`@      Z@     �d@     �b@      2@      @      .@      ,@               @      4@      �?      @      (@      1@       @      @              @      @                      @              �?      @               @       @      @      (@      @               @      *@      �?      @      "@      1@      @      @       @     �Y@     `c@      4@      4@      c@     �E@     @`@      W@     `b@     �a@      *@      �?      7@      O@              "@      J@      ,@     @Q@      B@     �O@     �I@      @      @     �S@     @W@      4@      &@     @Y@      =@     �N@      L@      U@     �V@      $@       @     �^@     pt@       @      7@      k@     �@@     ��@     �T@     8�@     �b@      @              9@     @X@              @     �B@      @     pu@      @     @g@      ;@       @              ,@     @P@              @      ;@      @     �g@       @     �R@      &@                       @      A@              @      4@       @     �[@       @      ?@       @                      @      ?@                      @      �?      T@              F@      @                      &@      @@                      $@      @      c@      @     �[@      0@       @              &@      @@                       @              b@             �V@      "@      �?                                               @      @       @      @      4@      @      �?       @     �X@     �l@       @      1@     `f@      ;@     �{@     @S@     �v@      _@      @              <@      S@       @       @     �P@       @     �V@      H@     �P@      ;@                       @      @              @      @       @              @      @      @                      :@     @Q@       @      �?      O@      @     �V@      F@      P@      6@               @     �Q@     @c@      @      "@     @\@      3@     @v@      =@     �r@     @X@      @       @      O@     �b@      @      "@     �Y@      1@     �u@      <@     �r@     @X@      @               @      @       @              &@       @      @      �?       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ%:hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @ĝA��R@�	           ��@       	                    @��JB�@�           ��@                          �5@��I?�@Q           �@                           �?���;M@�           ��@������������������������       �)�$�@�            �k@������������������������       ��aZ�Y;@           p{@                          �<@Nj�	�	@�           ��@������������������������       ��{1�q	@^           (�@������������������������       �� ���@S            �a@
                          �4@�����8@�            �@                           @Y�Y7�@�           ��@������������������������       �p���@r             g@������������������������       ��6`@�           8�@                           @2��� @�           H�@������������������������       ����\1p@           �z@������������������������       ��.8��@�            @k@                           @�`�5�@�           ��@                           �?�j����@           Њ@                           �?<9�C�@�            �k@������������������������       �g� @$             O@������������������������       ��Ot�@n             d@                           �?o�zװ	@�           ؃@������������������������       �T/	f��	@5           p@������������������������       �Q�B��@S            �`@                           �?��+7��@�            0r@                          �3@ҳԇ�?8            �X@������������������������       ��l#���?             J@������������������������       �'�֞� @             G@                           @w=�U¯@q             h@������������������������       ��zd΀ @<            �X@������������������������       �#j����@5            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `r@     �@      @@      H@     �{@     @Y@     ȏ@     �h@     H�@      u@     �B@      $@     �i@     0z@      ,@      <@     0q@     @S@     `�@     �a@     ��@     @l@      8@      "@     �_@      j@      "@      4@     �d@      J@     @m@      [@      p@      a@      5@      �?     �F@     @V@      @      @      S@      2@     `c@     �F@     �b@     �N@       @              0@      5@                      0@      @      O@      "@     �R@      .@              �?      =@      Q@      @      @      N@      (@     @W@      B@      S@      G@       @       @     �T@     �]@      @      *@     @V@      A@     �S@     �O@     �Z@      S@      *@       @     �P@      Z@      @      $@     �Q@      8@     �Q@     �F@     �V@      E@      *@              0@      .@              @      2@      $@      "@      2@      1@      A@              �?     �S@     `j@      @       @     �[@      9@     �@     �@@     0u@     @V@      @             �A@     �Z@      @      @     �@@       @     u@      @      h@      G@       @              *@     �D@                       @       @     �P@      �?      @@      4@                      6@     @P@      @      @      9@             �p@      @      d@      :@       @      �?     �E@     @Z@       @      @     @S@      7@      f@      ;@     @b@     �E@      �?      �?      >@     �P@       @      @      K@      "@      a@      (@     @V@      :@                      *@      C@                      7@      ,@      D@      .@     �L@      1@      �?      $@     @V@     @c@      2@      4@     @e@      8@     �p@      M@     �j@      \@      *@      $@     �S@      `@      ,@      1@     �b@      7@     �c@      L@     �^@     @V@      (@              0@      @@       @      �?      A@              S@      &@     �A@      0@                      @      $@                      @              @@       @      $@                              (@      6@       @      �?      >@              F@      "@      9@      0@              $@     �O@      X@      (@      0@     @]@      7@      T@     �F@      V@     @R@      (@      $@      K@      R@      &@      ,@      Y@      4@     �F@      <@     �S@      M@      (@              "@      8@      �?       @      1@      @     �A@      1@      "@      .@                      $@      :@      @      @      3@      �?     @\@       @     @V@      7@      �?              @      @               @      @              H@              @@       @                      @       @                                      8@              6@                               @      @               @      @              8@              $@       @                      @      5@      @      �?      0@      �?     @P@       @     �L@      5@      �?               @      @                       @      �?     �G@      �?      <@      @      �?               @      ,@      @      �?       @              2@      �?      =@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�#�ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���O@�	           ��@       	                   �2@�XƲ	�@~           t�@                           @\q���@2           @                           �?���ԕ@�             x@������������������������       �t����:@�             o@������������������������       ��B�2S@S             a@                          �0@��s��@@            �[@������������������������       �X|�P8Y�?             0@������������������������       ��[�i�@5            �W@
                           �?[%��B	@L           $�@                          �<@�*G���@8           P~@������������������������       �ix�pM@           �z@������������������������       �`C�@'            �N@                          �<@�u+7E�	@           ��@������������������������       �2��O`�	@�           x�@������������������������       �O�2b}@u            �h@                            @���F�g@/           <�@                           �?�y]�D�@{           �@                            �?;^�ڂ�@0           �~@������������������������       �����B@M            @_@������������������������       ��d��C@�            �v@                          �7@��hI�@K           x�@������������������������       ��P�Ȝ�@�           x�@������������������������       �w �[�]@�             l@                           �?ǔ[%Y@�            Pq@                          �4@���_q�?A            �Y@������������������������       ��<ę��?%             K@������������������������       ��x�b���?            �H@                           @LQ��2�@s            �e@������������������������       �Zܬ�M�@2            �Q@������������������������       � ��]@A            �Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     `@     �@@     �J@     `{@     @W@     (�@      l@     ؉@     �x@      4@      *@     @l@     `r@      5@     �C@     `r@     �P@     �x@     �g@     �x@     pq@      1@       @     �A@      R@      �?       @      H@      @     �b@     �A@      Y@      H@                      8@      H@      �?      �?      F@             @_@      4@      V@     �A@                      5@      =@      �?      �?      A@              P@      ,@     @P@      4@                      @      3@                      $@             �N@      @      7@      .@               @      &@      8@              �?      @      @      7@      .@      (@      *@                              @                      �?               @                                       @      &@      1@              �?      @      @      .@      .@      (@      *@              &@     �g@     �k@      4@     �B@     �n@      N@      o@     `c@     �r@     �l@      1@             �E@      S@      �?      @      O@      @     @X@      A@      [@      J@      @              D@     �Q@      �?      @      I@      @     �W@      8@     �Y@      A@       @              @      @               @      (@              @      $@      @      2@      �?      &@     �b@     @b@      3@      @@      g@      L@      c@     @^@     �g@     `f@      ,@      @     �^@      `@      2@      ;@      e@      F@      `@     @X@     �e@     �_@      ,@      @      :@      1@      �?      @      .@      (@      8@      8@      2@      J@               @     �V@      j@      (@      ,@      b@      ;@     ��@     �A@     �z@     �\@      @       @      U@      g@      @      "@     �^@      7@     P~@      @@     @v@     �W@       @              1@     �N@      �?      �?      ?@      @     �m@      "@     �[@      1@      �?                      (@      �?              (@       @      M@       @      >@       @                      1@     �H@              �?      3@      @     `f@      @      T@      "@      �?       @     �P@      _@      @       @     �V@      1@      o@      7@     �n@     �S@      �?             �G@      Y@      @      @     �L@      *@      k@       @      g@      J@      �?       @      4@      8@      �?      @      A@      @      ?@      .@      O@      :@                      @      7@      @      @      6@      @     �\@      @     @R@      3@      �?              @      @                       @             �N@      �?      =@      �?                       @      @                                      ;@              3@      �?                      �?      �?                       @              A@      �?      $@                              @      1@      @      @      4@      @      K@       @      F@      2@      �?              �?      @               @      .@      �?      ;@       @      &@      @                      @      $@      @      @      @      @      ;@             �@@      *@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�{dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @����E@�	           ��@       	                    @t['�@�           �@                           �?d���yh@T           ��@                           �?���W�@=           �@������������������������       ��v�*O@�            q@������������������������       �bB��=	@�           ��@                           �?o����@           �z@������������������������       ��&�7@|            �f@������������������������       ��(�y�e@�             o@
                           �?"/@��@�           H�@                            �?�5��	@:           X�@������������������������       �A�����?S            �`@������������������������       �_'(jC@�            @x@                           �?H-�6�@d           8�@������������������������       �wF��ҁ@#           0}@������������������������       �� �%E@A           @@                           @���@�            �@                          �3@p�%��@           ��@                          �1@�;'m3@�            @q@������������������������       �y���/�@C            �W@������������������������       �%'�$��@t            �f@                           @np��&	@`           �@������������������������       ��A�Ê-	@:           �}@������������������������       �3�Δ�7@&            �P@                           @����@�            pq@                           @��:�� @e            �d@������������������������       �7#��?O            �_@������������������������       ��#Q/eP�?             C@                           �?n�|$�@O            �\@������������������������       �OP`}1 @"             I@������������������������       ���8�B@-            @P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �q@     ��@      =@     �L@     }@      O@     ��@     �k@     �@     �u@      ;@      @     �k@     �w@      .@     �@@     �s@     �D@     ��@      b@     ��@     �n@      5@      @     �a@      f@      "@      4@     `g@      <@     �m@     �\@     �l@     @d@      1@      @      Z@     �_@       @      0@     @a@      3@     @`@     �T@     �`@     �]@      .@      �?      7@     �G@                      >@       @      K@      .@     �Q@      9@      @      @     @T@      T@       @      0@      [@      1@      S@      Q@      P@     @W@      $@             �B@     �H@      �?      @     �H@      "@     �Z@      @@      X@      F@       @              $@      8@               @      5@      @     �D@      3@     �B@      6@      �?              ;@      9@      �?       @      <@      @     �P@      *@     �M@      6@      �?      �?     �S@      i@      @      *@     @`@      *@     X�@      >@     pw@      U@      @              4@     @R@      @       @      B@      @     �o@      "@      Y@      4@       @                      ,@      @              $@      @     �R@      �?      9@      @                      4@     �M@               @      :@      �?     @f@       @     �R@      1@       @      �?     �M@     �_@      @      &@     �W@       @     �r@      5@     0q@      P@       @      �?      D@      O@       @      @      K@      @     �`@      $@     @]@      C@      �?              3@     @P@      �?      @      D@      @     @e@      &@     �c@      :@      �?      $@     �P@     �d@      ,@      8@     �b@      5@     �p@      S@     �h@     @Y@      @      $@     �M@     �a@      *@      4@     �_@      4@     �c@     @R@      [@      U@      @      @      *@     �F@      �?      @     �B@      @     �S@      (@      D@      =@                      @      ,@      �?      �?      $@             �B@      @      .@      @              @       @      ?@              @      ;@      @      E@      @      9@      7@              @      G@     �W@      (@      ,@     �V@      *@     �S@     �N@      Q@     �K@      @      �?      D@      S@      (@      ,@     @S@      (@     �Q@      I@     �P@      I@      @       @      @      3@                      *@      �?      @      &@      �?      @      �?               @      :@      �?      @      5@      �?     �[@      @      V@      1@                      @      .@                      &@      �?      Q@      �?     �M@      @                      @      .@                      @      �?     �L@      �?      E@                              @                              @              &@              1@      @                       @      &@      �?      @      $@              E@       @      =@      ,@                       @                      �?      @              7@       @      ,@      �?                              &@      �?      @      @              3@              .@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��rmhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?v,/�?G@�	           ��@       	                    �?��9��2	@	           l�@                           �?�DW�@A           x�@                          �1@�xK8x@|            �g@������������������������       ����#}W�?            �@@������������������������       ��ym���@g            �c@                           �?JjS;�@�             u@������������������������       ����qC�@b            `e@������������������������       ���S�@c            �d@
                           �?-{%�?�	@�           0�@                            �?����^@           �y@������������������������       ��b\��@K             _@������������������������       ��G�-u�@�            �q@                           �?�?��
@�           ��@������������������������       �,�9�	@�            �l@������������������������       ��.�W��	@&           �|@                          �4@\i�>�@�           ܡ@                           �?���"�@           (�@                          �0@I�L�= @            {@������������������������       ���b���?&            �M@������������������������       �#J��F# @�            pw@                           �?(�}��@�           ��@������������������������       �u�![�@            �F@������������������������       � ��k�@�           X�@                           @M `S@�           ��@                           �?�^$5��@U           (�@������������������������       ���١��@�            `s@������������������������       ��~nP�G@�           x�@                           �?f�=1��	@D            �W@������������������������       �J�!@             @@������������������������       ����hG	@,            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �t@     �@     �@@     �D@     p|@      V@     �@     �j@     ��@      v@      :@      3@      g@      n@      5@      8@     `n@     �J@     �i@      a@     �p@     �j@      5@       @      L@     �T@      @      $@     �R@      �?     @Y@      6@     �Z@     �P@       @       @      1@      7@                      =@             �K@       @     �F@      2@                      �?       @                      $@              .@              @      �?               @      0@      5@                      3@              D@       @     �D@      1@                     �C@      N@      @      $@     �F@      �?      G@      4@     �N@     �H@       @              1@      A@      @      @      4@      �?      9@      $@      <@      :@                      6@      :@              @      9@              5@      $@     �@@      7@       @      1@      `@     �c@      2@      ,@      e@      J@     �Z@     �\@     �c@     @b@      3@      �?     �B@      R@       @      @     �L@      ,@     �L@      B@     �L@     �P@      @              .@      *@              @      0@      @      6@      .@      6@      (@              �?      6@     �M@       @      @     �D@       @     �A@      5@     �A@     �K@      @      0@     �V@     @U@      0@       @      \@      C@     �H@     �S@     �Y@     �S@      0@      @      =@      G@      @      @      8@      0@      (@      <@      :@     �@@      @      (@      O@     �C@      "@      @      V@      6@     �B@     �I@      S@      G@      *@      �?      b@     �r@      (@      1@     �j@     �A@     ��@      S@     X�@     �a@      @              M@     �d@      @      $@     �S@      @     0�@      A@     r@      N@       @              6@      G@              @      2@             �l@      @     @X@      ,@       @                      1@                       @              <@              $@       @                      6@      =@              @      0@              i@      @     �U@      (@       @              B@     @^@      @      @      N@      @      r@      >@      h@      G@                      @      @              �?      &@      �?      (@      �?      @      @                      @@     �\@      @      @     �H@       @     `q@      =@     @g@     �E@              �?     �U@     �`@      @      @     �`@      @@     �p@      E@     �p@     @T@      @      �?     �R@     �^@      �?      @     �]@      =@      p@      ?@     �o@      R@                      3@     �B@                      ;@       @     @]@      @     �R@      5@              �?      L@     @U@      �?      @      W@      5@     `a@      9@     @f@     �I@                      (@      (@      @      �?      .@      @      (@      &@      *@      "@      @              @      @              �?       @               @      @      @               @              @      "@      @              @      @      $@      @      @      "@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�v��0@�	           ��@       	                    �?p�&�@j           �@                          �:@�òy6	@�           ��@                           �?�^O�@           x�@������������������������       ��.}��:@4           �@������������������������       ���ۇ1	@�           0�@                           �?L,PU��	@�            �t@������������������������       ��B��Z@@            �Y@������������������������       � 

@�             m@
                          �1@�5H.�@           ��@                            @����g@6             W@������������������������       �2��>C@%             M@������������������������       ����IEQ�?             A@                          �4@�/��5*@I           �@������������������������       �g���@�             j@������������������������       �ava|�I@�            �r@                          �1@���@G           �@                           @:�O( @�             w@                           @US).��?}             h@������������������������       �6�<B��?G            �]@������������������������       �R�]E@6            �R@                           @�4���@s             f@������������������������       ���]]ȍ @F             [@������������������������       ��V��q5@-            @Q@                           �?��ќU�@W           P�@                           �?� ���@           �z@������������������������       �H�q��o@�            �m@������������������������       �- |�}�@r            �g@                          �<@��q��q@U           P�@������������������������       ���+J?@0           Ћ@������������������������       �?p�GM @%             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     `q@     ��@      9@     �K@     �~@      W@     ��@     `h@     ��@     w@      5@      5@      i@     @t@      0@      E@     Pu@      R@      w@     �d@     �v@      o@      3@      5@      d@     �l@      .@      C@     �p@      J@     `l@      ]@     @n@     �h@      3@      @     �^@     @i@       @      @@     �i@     �@@     �h@     �T@     `j@     �_@      0@       @      <@     @T@      �?      "@      U@      "@     @\@      >@     @V@     �K@      @      @     �W@     @^@      @      7@     �^@      8@     @U@     �J@     �^@      R@      *@      ,@     �B@      :@      @      @     �N@      3@      =@     �@@      ?@     @Q@      @       @      @      @      @              <@      @      (@       @      @      :@       @      (@      >@      4@      @      @     �@@      0@      1@      9@      9@     �E@      �?              D@      X@      �?      @     �R@      4@     �a@      H@     �^@      J@                       @      2@                      @              C@      &@      3@      �?                       @      @                      @              9@       @      *@                                      &@                                      *@      @      @      �?                      C@     �S@      �?      @     �Q@      4@     �Y@     �B@     �Y@     �I@                      $@      ?@      �?       @      F@      @      A@      "@      J@      6@                      <@     �G@               @      ;@      1@     @Q@      <@     �I@      =@              �?     �S@     �m@      "@      *@     `b@      4@     (�@      ?@     �z@     @^@       @               @      A@              @      7@             �h@      @     �U@      *@      �?              @      *@              �?      @             �_@      �?      A@      @      �?              @      @                      �?             �V@              1@       @                       @      "@              �?      @              B@      �?      1@       @      �?              �?      5@              @      1@             �Q@      @      J@      "@                      �?      &@                      ,@             �A@             �D@      @                              $@              @      @             �A@      @      &@      @              �?     �Q@     �i@      "@       @      _@      4@     |@      ;@     `u@      [@      �?              0@      M@      �?      �?      9@      @     �g@       @     �Y@      4@                      &@      9@              �?      0@      @     @^@      @      G@      &@                      @     �@@      �?              "@             @Q@      @     �L@      "@              �?      K@     `b@       @      @     �X@      0@     0p@      3@     �m@      V@      �?      �?     �I@     �a@      @      @     @U@      0@      p@      2@     �l@     �S@      �?              @      @       @              ,@              @      �?      $@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJfG�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��u�/@�	           ��@       	                    �?!�+���@�           �@                          �<@+�)B��@�           ��@                          �3@��qe�@p           x�@������������������������       ���s�:�@�             n@������������������������       ��Nt��@�            �s@                            �?�&[06@+            �P@������������������������       ��Qlc$@            �C@������������������������       ���2h�.@             ;@
                           �?0̾�=	@�           p�@                           �?6{�Hn�	@�           Б@������������������������       �Ӌ �	@�             x@������������������������       �}Hu�	@�           ��@                           �?��P,y�@           �z@������������������������       ����ڵ@             @@������������������������       �d� �1�@�            �x@                          �4@PQt�S@1           �@                           @�G��@R            �@                           �?8Yt˥\@�            �j@������������������������       �f�n�@J            @[@������������������������       �By!��@J            @Z@                            �?Z�J�
@�           p�@������������������������       �����{g@�             y@������������������������       ��[0-�+ @�            �s@                           @G�K�p�@�           ��@                          �5@,�]N�@0           `@������������������������       �e�-�7�@@            �]@������������������������       ���ʁ�@�            �w@                           @zċ��@�             r@������������������������       ����=ɤ@`            �c@������������������������       ��H���U@O            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@      �@      9@      P@     �z@     �S@     �@     @i@     �@     �u@      =@      .@      l@     0t@      4@     �F@     �q@     �N@     �w@      e@     �x@     `o@      7@      �?     �N@      Q@       @      @     @P@      @     �d@      C@     �b@      L@      @      �?      L@      N@       @      @      L@      @     �d@      >@     �`@     �C@      @              ,@      6@                      5@              T@      *@      P@      :@              �?      E@      C@       @      @     �A@      @     @U@      1@     �Q@      *@      @              @       @              @      "@              �?       @      ,@      1@      �?               @      @                      @                       @       @      ,@      �?              @      @              @      @              �?              @      @              ,@     `d@     �o@      2@      C@     @k@     �K@     �j@     @`@     �n@     `h@      1@      ,@     �`@     �e@      .@      =@      e@      F@     ``@     �V@      f@     `b@      1@      @     �E@     �R@      @      @      J@      ,@      H@      >@     �D@      N@       @      &@     @V@      Y@      $@      8@      ]@      >@     �T@     �N@      a@     �U@      "@              ?@      T@      @      "@      I@      &@      U@     �C@     @Q@      H@                      �?      @              "@       @      @      �?      @       @      @                      >@     �R@      @              H@       @     �T@      B@     �P@     �E@              �?     �W@     �o@      @      3@      b@      1@     H�@      A@      y@      Y@      @             �E@      _@      @      "@     �E@      @     �{@      *@     �i@     �F@      @              3@     �G@                      &@      @     �S@      @      D@      (@                      0@      8@                       @              B@      @      0@      @                      @      7@                      @      @      E@              8@      @                      8@     @S@      @      "@      @@             �v@      $@     �d@     �@@      @              &@      G@      @      @      7@              g@      @     �Y@      5@                      *@      ?@              @      "@              f@      @     �O@      (@      @      �?     �I@      `@       @      $@     @Y@      *@      j@      5@     �h@     �K@      @      �?     �A@     �Q@               @     �P@      "@      d@      "@     �^@      7@      @              �?      ;@                      5@      �?      <@      �?     �A@       @      @      �?      A@     �E@               @      G@       @     �`@       @     �U@      5@                      0@     �M@       @       @      A@      @      H@      (@     �R@      @@                      �?     �E@       @      �?      *@      @     �@@      $@      D@      $@                      .@      0@              @      5@      �?      .@       @     �A@      6@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJQZ�&hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�{�IF@�	           ��@       	                   �1@����P@n           �@                          �0@wA�Tă@t            �@                           �?x�ܢ��@y            �i@������������������������       ��<�R�?:             Z@������������������������       �{�3�@?             Y@                           �?Wh��0}@�            �w@������������������������       �O��a'@z             f@������������������������       �\�f+t@�             i@
                           �?X��,�Q@�           ��@                           @���)�@�            0z@������������������������       �����v@�             l@������������������������       �����'��?y            @h@                           @�e��E@�           ��@������������������������       �g�Kwj@Z           ��@������������������������       �=a���@�             p@                           @�^�1�f@T           ��@                           �?"V��XL	@M           h�@                           �?��.`�y@�            v@������������������������       ���a@�            �p@������������������������       ���r�'@2            �U@                           @����w	@i           ȍ@������������������������       ����bM	@           ؉@������������������������       �=��N�@Q            �_@                          �7@��ʤ��@           `�@                          �5@��/Xn@	           �z@������������������������       ����2R@m             f@������������������������       ���d�h@�             o@                          @@@����[@�             x@������������������������       ��?�Y7@�             w@������������������������       �i	\��p @
             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     @t@     p�@      >@      K@     `}@     �U@     ��@     �f@     ��@     �v@      7@      @     @Z@     �l@      @      1@     �e@      1@     ��@     �O@      z@      c@      (@              5@     �P@              @     �G@             �o@      *@     �`@     �C@       @              @      :@              @      2@             �T@              I@      4@                              &@                      @             �I@              <@       @                      @      .@              @      (@              @@              6@      (@                      1@      D@              @      =@             @e@      *@     �T@      3@       @               @      0@              @      (@              U@      @      B@      (@                      "@      8@                      1@             �U@       @     �G@      @       @      @      U@     `d@      @      &@     �_@      1@     pu@      I@     �q@     �\@      $@              >@      N@              @      9@      @     �b@      *@     @\@      7@                      2@      D@               @      1@      @      F@      &@      Q@      6@                      (@      4@               @       @              Z@       @     �F@      �?              @      K@     �Y@      @      @     @Y@      ,@     `h@     �B@     �e@     �V@      $@       @      C@      S@      @      @     �R@      "@      `@      $@     �^@      Q@      �?      @      0@      ;@       @      �?      ;@      @     �P@      ;@     �H@      7@      "@      2@     `k@     �t@      7@     �B@     �r@     @Q@      x@     @]@     �x@     �j@      &@      1@     �c@     @j@      2@      =@     �j@      J@      d@      Y@     @h@      b@      $@      @      E@      J@       @      @      L@       @     @U@      2@      L@      :@      @      @      @@      F@       @      @     �G@      �?      G@      0@     �E@      7@      @              $@       @                      "@      �?     �C@       @      *@      @      �?      ,@     �\@     �c@      0@      6@     �c@      I@      S@     �T@     @a@     �]@      @       @      X@     �`@      0@      6@     �a@      D@     @P@     �O@      `@     @Z@      @      @      2@      7@                      .@      $@      &@      3@      "@      ,@      �?      �?     �O@     �]@      @       @     �T@      1@      l@      1@     �i@      Q@      �?              @@     �R@      @       @      G@      $@      a@       @     �X@      4@                      @      >@              �?      3@      "@      K@      �?     �J@      @                      <@     �F@      @      �?      ;@      �?     �T@      �?      G@      ,@              �?      ?@      F@      �?      @     �B@      @     @V@      .@     �Z@      H@      �?      �?      :@      F@      �?      @     �B@      @     @V@      *@      Y@      G@      �?              @                                      �?               @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJD`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?F�E��H@�	           ��@       	                    �?Υ6W	@�           ؘ@                          �4@���L�@�           @�@                           @8��z�@�            �o@������������������������       ��ծ�@P            @`@������������������������       �����@W            �^@                           @[��ro@�            �t@������������������������       �3�KpnA@�            �r@������������������������       �6��-@             ?@
                          �7@�V�ֺ�	@m           p�@                          �4@��x���@w           h�@������������������������       �Y�7�_@�            x@������������������������       ���˫��@�            �m@                           @�6o=�i
@�            x@������������������������       ��^���@�             m@������������������������       ��+�"@`             c@                           �?��8�64@�           &�@                           �??bEq�@�           (�@                           @x�anm'@�            y@������������������������       ��B�[@6            @V@������������������������       ���I�D�?�            �s@                           @M��pQ
@�            @u@������������������������       ��t� Vb@�            Pp@������������������������       � 9�y
�@8            �S@                          �4@Z�*��R@�           ��@                           @E���'@�           `�@������������������������       �3�R�V@|            @j@������������������������       �#2�R�a@n           Ё@                          �7@��j�@�           �@������������������������       ����}@�            0y@������������������������       �ܖO�@�            �x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     (�@      9@     �J@     �{@      R@     ��@     �n@     ��@     �v@      >@      0@      g@     �l@      4@      >@     @m@     �C@     �l@     �_@     @p@     `i@      5@      �?      G@      Y@       @       @     @V@      @     @Z@      D@     �Z@     @R@      @      �?      .@     �G@                      A@      �?     �I@      ,@      M@      ?@      �?      �?      @      :@                      0@              :@      @      E@      $@                      $@      5@                      2@      �?      9@      $@      0@      5@      �?              ?@     �J@       @       @     �K@      @      K@      :@      H@      E@      @              :@      J@       @       @     �G@      @     �J@      2@      H@     �A@      @              @      �?                       @              �?       @              @      �?      .@     @a@      `@      2@      6@      b@      @@     �^@     �U@     @c@     @`@      ,@      "@     @U@     �R@       @      &@     �V@      @     @X@      E@     �\@      S@      @      @      E@     �@@      @      $@      N@       @     �R@      =@     �Q@      I@      @      @     �E@      E@       @      �?      ?@      @      7@      *@      F@      :@              @     �J@     �J@      $@      &@      K@      9@      :@     �F@     �C@      K@      "@       @      @@      F@       @      @     �D@      "@      .@      1@      7@     �C@       @      @      5@      "@       @      @      *@      0@      &@      <@      0@      .@      @       @     @`@     t@      @      7@     �i@     �@@     ��@      ^@     x�@      d@      "@              :@     �U@      �?      @      E@      @     �u@      2@     `f@     �@@      @              (@      F@              @      ?@      �?     @j@      $@     �Q@      3@                      @       @              @      .@      �?     �A@      @      .@      @                      @      B@                      0@             �e@      @     �K@      0@                      ,@      E@      �?              &@      @     �`@       @     @[@      ,@      @              ,@      A@                      @      @      [@      @     @T@      "@       @                       @      �?              @              :@      @      <@      @       @       @      Z@     `m@      @      3@     �d@      =@     �{@     �Y@     �u@     �_@      @             �D@     �\@      @      @      J@      @     �r@     �H@     �d@      F@                      @      C@              @      3@      �?     �R@      A@      8@      (@                     �B@      S@      @      @     �@@      @     �k@      .@     �a@      @@               @     �O@     @^@      �?      *@      \@      7@      b@     �J@     �f@     �T@      @              =@     �N@      �?      @      M@      .@     �V@       @      Y@      ?@      @       @      A@      N@              "@      K@       @      K@     �F@     @T@      J@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��{ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��4Ufr@�	           ��@       	                   �4@:q{�\@"           4�@                           @g�bX�@h           �@                           @-����@h            �@������������������������       ���]~a @�            0v@������������������������       �)^=*�1@|             h@                           �?�wHR@            �@������������������������       �F�pl�Y�?�            @q@������������������������       ��D�(��@K           H�@
                           �?�-��p@�           d�@                           @;��>�	@�           ��@������������������������       ���+V	@X           ��@������������������������       �Z3�4�	@4             U@                           @Fĥ�$�@.           H�@������������������������       ��l��^2@�            �w@������������������������       ���lf@=           �~@                           �?��P9Q@�           ��@                          �<@�z#��i	@�            �@                          �1@?aAGJ7	@c           p�@������������������������       ��?j�n=@'            �N@������������������������       ��rN��\	@<           @                           �?��h�@1            �T@������������������������       ��/ѕ��@            �C@������������������������       � %[��@            �E@                          �3@��oT�@           �z@                           @ �&�'@r            `g@������������������������       �o�Ӱd@-             S@������������������������       �+?�F���?E            �[@                           @Q��bL)@�            �n@������������������������       ��؇�?@<            �V@������������������������       ��v*8B�@f             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     ��@     �@@     �L@     P}@     �U@     X�@      m@     Ȉ@     �u@      B@      @     �j@     �x@      4@     �C@     �s@     �L@     ��@     @e@     ��@      o@      5@      �?      P@      g@      @      @      ]@      $@     0~@     �T@     r@     �X@      @      �?      9@     @U@      @      @     @Q@      @      `@     �P@     �Y@     �K@      @              3@     �G@              @     �E@      �?     @V@      >@     �S@      E@      �?      �?      @      C@      @      �?      :@      @      D@      B@      8@      *@       @             �C@      Y@      @       @     �G@      @      v@      1@     @g@     �E@                      .@      >@                      @             @d@      @     �I@       @                      8@     �Q@      @       @     �D@      @      h@      *@     �`@     �A@              @     �b@     �j@      ,@      @@     @i@     �G@     0q@     �U@      s@     �b@      2@      @     �O@     �V@      "@      1@     �Z@      5@     �Q@     �J@     @X@      S@      ,@      @     �M@     �T@       @      1@      V@      *@     �P@      B@     @W@      Q@      @      @      @      @      �?              3@       @      @      1@      @       @       @             @U@     �^@      @      .@     �W@      :@     �i@      A@      j@     �R@      @              E@     �E@               @     �C@      3@      Y@      2@     @R@     �B@      �?             �E@     �S@      @      @      L@      @      Z@      0@      a@     �B@      @      @     @Y@     �`@      *@      2@     �b@      >@     �n@     �O@     �h@     �X@      .@      @     �S@     �U@      (@      "@     �Z@      4@      T@      I@     �Y@      S@      *@      @      P@      Q@       @      @      W@      3@     �S@     �E@     �W@     �P@      *@              @      @       @              @              3@      �?      $@      $@              @      M@      O@      @      @     @U@      3@      N@      E@     @U@      L@      *@       @      .@      2@      @      @      ,@      �?      �?      @      @      $@               @      �?      *@       @              (@      �?      �?      �?      @      @                      ,@      @       @      @       @                      @      @      @                      6@      G@      �?      "@     �F@      $@     �d@      *@      X@      6@       @              @      2@              @      @             �V@      @     �G@      @                              *@              @                      ?@      @      .@      @                      @      @                      @              N@              @@      �?                      .@      <@      �?       @     �C@      $@     �R@       @     �H@      0@       @               @      1@                      2@      @      6@      @      $@      @                      @      &@      �?       @      5@      @      J@      �?     �C@      (@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�͈hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @yu��Xo@�	           ��@       	                    �?�J��8 @�           Υ@                           �?p!X@H           p�@                           �?h���Z�@?           h�@������������������������       ��;�@Z             c@������������������������       �۽�C38@�            Pw@                           @��E�·@	           z@������������������������       ����@�            `m@������������������������       �8�Q��|@t            �f@
                          �4@�[��@�           �@                          �1@6��ʟ>@�           ��@������������������������       �-A-� @�            �o@������������������������       �w���@Z           ��@                           @�@D�C	@�           t�@������������������������       ���$�	@�           ��@������������������������       ��ܦE��@           `|@                           �?�xL�J@�           ��@                          �8@��_f	@�           P�@                           @�Z<�Jd@/            }@������������������������       ��	��R@�            �r@������������������������       �������@m            `d@                           �?��)�
@�            @k@������������������������       �z(3O�(@             J@������������������������       �h$8�	@a            �d@                           �?�':��@           �{@                           @9�Fr�@�            @k@������������������������       ����J@>            �U@������������������������       ����W@P            �`@                           @f�0�*/@�            �k@������������������������       �����A@<             X@������������������������       ��3��w@S            �_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pt@     x�@     �D@     �I@     �{@     @S@     P�@     �l@     ��@     �u@      @@      "@     �j@     py@      3@      >@     `r@      L@     ��@     �e@     ��@     �n@      4@             �Q@     @`@               @     @T@      $@     �u@     �A@     `h@     @P@      @             �B@      W@               @     �F@      "@     `i@      6@     �S@     �A@       @              2@      B@              �?      0@      @      @@      2@      "@      0@       @              3@      L@              �?      =@      @     `e@      @     @Q@      3@                     �@@      C@                      B@      �?     `b@      *@     @]@      >@       @              :@      3@                      ;@             �L@      @      T@      2@       @              @      3@                      "@      �?     �V@      @     �B@      (@              "@     �a@     Pq@      3@      <@     �j@      G@     �y@     @a@     @w@     �f@      0@      �?      E@     �Z@      @      @     @R@      @      o@      I@     `g@     �R@       @      �?      @      >@                      1@      �?     �W@      ,@     �P@      7@                     �B@      S@      @      @      L@      @     @c@      B@      ^@      J@       @       @      Y@     `e@      .@      9@     �a@      E@     �c@      V@      g@     �Z@      ,@      @     @Q@     @W@      "@      3@      S@      >@      Q@      Q@      V@     @P@       @       @      ?@     �S@      @      @      P@      (@     �V@      4@     @X@     �D@      @      "@     @\@      c@      6@      5@     �b@      5@     �n@      L@     @k@     @Z@      (@      "@     �T@     �X@      1@      *@     @\@      0@      V@     �F@     @\@     �R@      (@       @      F@     �O@      @       @     �V@      @     �R@      6@     �U@     �I@      @      @      @@      E@      @       @     �L@      @     �P@      $@     �J@      9@      �?      @      (@      5@              @     �@@      @       @      (@     �@@      :@      @      �?      C@      B@      (@      @      7@      $@      ,@      7@      ;@      8@      @              ,@      @      �?              @       @      @              @      @      @      �?      8@      >@      &@      @      0@       @      @      7@      5@      2@       @              ?@     �J@      @       @      B@      @     �c@      &@     @Z@      >@                      $@      1@      @      �?      *@      @     @V@      @      M@      0@                      @      (@      �?              @       @      =@      @      2@      @                      @      @      @      �?      @      @      N@              D@      "@                      5@      B@              @      7@             �P@      @     �G@      ,@                      &@      ;@              @      @              ?@      @      "@      @                      $@      "@              @      1@              B@      @      C@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJx"�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��~1U@�	           ��@       	                   �5@O�F��@^           �@                          �1@q��.��@�           ��@                           @H�#���@�            �o@������������������������       ���
+�@�            �m@������������������������       ��"��~@
             3@                           �?K���;@
           �@������������������������       ��n��y@�            �o@������������������������       ��2n�	@k            �@
                          �;@ȸ��5�	@�           ��@                          �7@�lؽ��@�           ��@������������������������       �~�h��@�            `u@������������������������       � g�6	@*           �}@                           �?o7�,�	@�            Ps@������������������������       �<��?'C@6            @V@������������������������       �ZLi��
@�            �k@                            @��?�@1           ��@                           @�@��8�@�           p�@                          �5@��(�t@�           X�@������������������������       ���ܟ��@�           H�@������������������������       �S%d�@@�            �t@                           �?�8#��@�            `x@������������������������       �$���K
@a            `c@������������������������       �uH98ɲ@�            `m@                          �9@^�Ր�@�             r@                          �5@����8@�             o@������������������������       ��8jS/� @l             g@������������������������       ��sr��"@'             P@                           @b�K���@             E@������������������������       ��	�U$	�?             3@������������������������       �aA�6�@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     ��@      9@      N@      }@     �T@     (�@     �m@     ��@     @w@      ?@      ,@     �h@     `r@      3@      G@     pt@     �Q@     `v@     @h@      x@     �o@      =@      @      O@     �a@      @      9@     �b@      5@     �m@     @S@     �k@     �Z@       @              "@     �B@               @      F@              Q@      ,@      L@      9@                      @     �B@               @     �B@             �P@      ,@      J@      6@                      @                              @               @              @      @              @     �J@     �Y@      @      7@      Z@      5@     @e@     �O@     �d@     @T@       @              2@      =@      �?      @      6@       @      T@      0@      P@      1@      �?      @     �A@     �R@      @      3@     �T@      3@     �V@     �G@     �Y@      P@      @      &@      a@     @c@      (@      5@     `f@     �H@      ^@     @]@     @d@     �b@      5@      �?     �Z@     �\@      @      *@     �`@      9@     �X@     �U@     �`@     �U@      3@      �?      O@      I@       @       @     �L@      @      A@      :@      K@     �E@      �?              F@      P@      @      @     @S@      5@     @P@      N@     �S@     �E@      2@      $@      >@      D@      @       @     �F@      8@      5@      ?@      >@      O@       @              &@      .@               @      *@              @      "@      .@      0@      �?      $@      3@      9@      @      @      @@      8@      ,@      6@      .@      G@      �?             @V@      o@      @      ,@      a@      (@     ��@     �F@     �y@     �]@       @             �T@     �k@      @      "@     �[@      &@      �@      E@     0u@     @Y@                      H@      d@      �?      @     �Q@      @     �y@      <@     �n@     �R@                      6@     �Z@              @      >@       @     �s@      0@     `f@     �D@                      :@     �J@      �?             �D@      @      X@      (@      Q@     �@@                      A@      O@       @      @      D@      @     �Z@      ,@      W@      ;@                      @      >@       @      �?      (@             �N@      @      @@      "@                      =@      @@              @      <@      @      G@      &@      N@      2@                      @      ;@      @      @      :@      �?     �^@      @      S@      1@       @              @      :@              �?      1@      �?     �Z@              R@      0@       @              @      1@              �?      ,@             @V@              H@      @       @                      "@                      @      �?      2@              8@      "@                      �?      �?      @      @      "@              0@      @      @      �?                                                       @              *@              @                              �?      �?      @      @      @              @      @              �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�œhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�L
�W@�	           ��@       	                    �?��E���@�           ��@                           �?��	#3@�           0�@                          �<@���l�@A           �@������������������������       �m�ճ1@           0|@������������������������       �H�1��@&             N@                          �<@^}oCL@q            �d@������������������������       �2q�c�@j            �c@������������������������       ��tc��@             &@
                          �9@,���c	@�           ��@                           �?fY+��@�           t�@������������������������       ����q�T	@           0�@������������������������       ���{�K0@�            pu@                           �?���x	@�            y@������������������������       �cg�%_"@O            �a@������������������������       �&T|��*	@�            Pp@                           @T�ݾ��@%           ԙ@                            �?�=���@�           �@                           @r���v�@�           ��@������������������������       �'..��@�            @k@������������������������       ������@�            Px@                          �3@�>��@S            �@������������������������       �R��P� @�            `o@������������������������       ��"R���@�            �r@                           �?���]T@G            @                          �3@��e�@�            �m@������������������������       ����	�G@;            �W@������������������������       ����&�a@d            �a@                           @�#Z�/@�            `p@������������������������       �l""�>�@M            �`@������������������������       ��/\r�@[            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pt@     �@      9@      I@     P~@     �Q@      �@     �m@     ؉@     w@      ?@      3@     �n@     �s@      3@     �D@      u@     �M@     0w@      i@     �w@     `o@      8@       @     �V@     @U@              "@     �R@      @     `e@      ?@     �b@      N@       @       @     �Q@     @R@              "@     �L@       @      \@      <@     �Z@     �H@       @       @      P@     @P@              @      H@       @     �[@      8@     �X@      >@       @              @       @              @      "@              �?      @      @      3@                      3@      (@                      1@      �?     �M@      @     �F@      &@                      .@      (@                      0@      �?      M@      �?     �E@      $@                      @                              �?              �?       @       @      �?              1@     `c@     �l@      3@      @@     �p@      L@      i@     @e@     �l@     �g@      6@      @     @]@     �f@      *@      >@     @i@      =@      f@     �[@     `f@      ^@      0@      @     �X@      `@      *@      7@      b@      4@     @X@      T@      ^@      W@      ,@              2@     �J@              @     �L@      "@     �S@      ?@     �M@      <@       @      &@      C@      G@      @       @      O@      ;@      8@     �M@     �H@     �Q@      @      @      "@      3@      @      �?      A@      (@              4@      "@      8@       @      @      =@      ;@       @      �?      <@      .@      8@     �C@      D@     �G@      @              T@     @i@      @      "@     `b@      (@     h�@     �A@      |@     �]@      @             �K@      `@      �?      @     @X@      @      }@      9@     �r@     �P@      @              9@      P@      �?              C@      @     �n@      2@     �d@     �F@       @              @      ?@                      $@      @     �U@      @      E@      <@       @              2@     �@@      �?              <@      �?     �c@      &@     �^@      1@                      >@     @P@              @     �M@      �?     �k@      @      a@      6@      @              $@      D@              �?      *@      �?     �\@      @     �P@       @                      4@      9@               @      G@              [@      @     �Q@      4@      @              9@     @R@      @      @      I@      @     �^@      $@     �b@     �I@       @              *@     �E@              @      7@      �?     �M@      @     �O@      9@                      "@      .@                      $@              ?@              ;@      @                      @      <@              @      *@      �?      <@      @      B@      6@                      (@      >@      @              ;@      @      P@      @     @U@      :@       @               @      3@      @              $@      @      9@      @     �G@      *@       @              $@      &@      �?              1@             �C@      �?      C@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJTu|hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�<g��W@�	           ��@       	                    �?�l$� 	@a           ��@                          �<@�����@�           ��@                           �?�~�� �@y           ��@������������������������       �i�Gs��@�            �q@������������������������       ��N�E�@�            �s@                          �?@t{�Y@2             W@������������������������       �����@$            �P@������������������������       �����@             :@
                           �?Fl��	@�           (�@                           �?�G�t.8	@G             ]@������������������������       ��%~@             A@������������������������       ��I��<�@0            �T@                           @[����l	@o           X�@������������������������       �1���2	@�           (�@������������������������       �*���	@�            �i@                           �?�_�@9           <�@                          �4@䏼�/U@r           ؂@                           @�+*�q�?�            �w@������������������������       ���*���?            �h@������������������������       �@Ⱦ%@h            �f@                           �?�<���`@�             l@������������������������       �q���@P            @`@������������������������       ��	��5�@;            �W@                          �1@NB���@�           Б@                           @o���	8�?u             f@������������������������       ���yEY�?P             ^@������������������������       ��ˏ�`-�?%             L@                           !@:ݱ�@R            �@������������������������       �m�|u�r@K           ��@������������������������       ����� � @             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      <@     �H@      |@     �S@     <�@      n@     @�@     Pv@     �C@      3@     �i@      s@      9@      B@     t@     �N@     @x@      h@     �u@     �m@     �A@              R@     @V@      �?       @     �T@      @     �e@     �E@     ``@      S@      @             �O@     �R@      �?       @     �P@      @     �e@     �B@      _@      H@       @             �@@      =@      �?      �?      C@      @     �S@      8@      J@      6@      �?              >@     �F@              �?      <@       @     �W@      *@      R@      :@      �?              "@      .@              @      0@              @      @      @      <@       @               @      ,@              �?       @               @      @      @      ;@       @              @      �?              @       @              �?       @      �?      �?              3@     �`@     �j@      8@      <@     �m@      K@     �j@     �b@     �j@      d@      ?@      @      "@      .@              @      :@      @       @      4@      "@      *@      @      �?       @      *@                      @       @              @      �?      @              @      @       @              @      3@      �?       @      0@       @      "@      @      *@     @_@      i@      8@      5@     �j@     �I@     `j@      `@     �i@     �b@      9@      $@     @Z@     �e@      8@      3@     �f@     �A@      g@      X@     �g@      `@      1@      @      4@      ;@               @      >@      0@      ;@     �@@      2@      4@       @      �?     �W@      m@      @      *@      `@      2@     X�@      H@     �z@      ^@      @              3@     @V@      �?      @      >@      @     �q@       @      a@      7@                      .@      D@              @      *@             �j@      @      T@      (@                      "@      4@                                      _@      �?      D@      @                      @      4@              @      *@             @V@       @      D@      @                      @     �H@      �?              1@      @     @R@      @     �L@      &@                      @      <@                      *@      @     �F@      @      ;@      @                              5@      �?              @      @      <@              >@      @              �?     �R@     �a@       @      $@     �X@      &@     �v@      D@     Pr@     @X@      @               @      ;@               @      @             @T@      �?      J@      @                       @      9@                      @             �F@              E@      @                               @               @       @              B@      �?      $@      @              �?     @R@      ]@       @       @     �W@      &@     �q@     �C@      n@     �V@      @      �?      R@     �\@       @       @     @W@      @     �q@     �C@     �m@     �V@      @              �?       @                      �?      @                      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�Z�i"`@�	           ��@       	                    @�7
DiX@�           ,�@                           �?�͹B�@J           ��@                           �?xs���@�            �q@������������������������       ��W6�a�@U            �_@������������������������       �ԥ���@c             d@                           @��\� l@�           ��@������������������������       ��0���'@�            �@������������������������       ��ȯ]"@             2@
                          �0@E��\�@I           ��@                           @/��{���?F            �\@������������������������       �<�8��\�?)            �P@������������������������       �ܿ=a5_�?            �H@                           �?n����$@            �@������������������������       ��QƤg��?�            �s@������������������������       �i����@J           `�@                           @ݐ�<�@           ��@                          �8@E2c�ɰ	@-           `�@                            @4X���@�           Є@������������������������       ��O��C	@�            �x@������������������������       ��m�e@�            �p@                           �?ٵ�ɭ�	@�           ��@������������������������       �ЉX���@j             e@������������������������       �w�\�M
@1           P}@                            @t���@�           0�@                            �?]l �7@�           ��@������������������������       ��� `��@�            `x@������������������������       �n��@�            �j@                           �?�|�N��@Y            @a@������������������������       ���R.��?             D@������������������������       ��;^��@?            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �q@     x�@     �@@      M@     �}@     �T@     ,�@     �k@     �@     �t@     �@@      @     �Z@      n@      "@      1@     �h@      2@     P�@     �W@     �x@     @_@      &@      @     �P@     �\@      @      &@      a@      0@      j@     @R@     �f@     �V@      "@              5@      @@               @      B@       @     @V@      .@     �Q@      1@      �?              @      &@              �?      6@       @      D@      (@      8@      @      �?              ,@      5@              �?      ,@             �H@      @     �G@      &@              @      G@     �T@      @      "@     @Y@      ,@     �]@      M@     �[@     @R@       @      @      E@     �T@      @      "@     �X@      ,@     �]@     �K@      [@     @R@      @      �?      @                              @              �?      @       @              @             �C@     �_@      @      @     �N@       @     �{@      6@     �j@     �A@       @               @      3@                      @             �O@              3@      "@                       @       @                      @             �C@              ,@                                      &@                                      8@              @      "@                     �B@     �Z@      @      @      M@       @     �w@      6@     @h@      :@       @              *@      5@              @      6@              f@      @     �N@      @       @              8@     �U@      @      @      B@       @     @i@      0@     �`@      3@              3@     `f@     �s@      8@     �D@     �q@     @P@     x@      `@     pw@      j@      6@      2@     �`@     �i@      2@     �A@     �h@      K@     `f@     @Z@     �g@     �b@      4@      "@     �S@     �Y@      @      7@     �Z@      8@      Z@     �@@      ]@     �L@      @      @     �I@      E@      @      3@     @P@      5@      P@      9@     �R@      7@       @      @      <@     �N@              @      E@      @      D@       @     �D@      A@      @      "@      L@     �Y@      (@      (@     @V@      >@     �R@      R@     @R@     @W@      .@              1@     �@@              @      :@      @      :@      @      9@      9@      @      "@     �C@     @Q@      (@       @     �O@      ;@     �H@     @P@      H@      Q@      (@      �?      F@     �\@      @      @      U@      &@     �i@      7@     @g@     �M@       @      �?     �B@     �Z@      @      @     �R@      &@      c@      6@      b@      G@       @              ;@     @R@       @      @     �A@       @     �X@      2@      X@      >@              �?      $@     �@@      @             �C@      @     �K@      @      H@      0@       @              @       @      �?      @      $@             �J@      �?      E@      *@                      @      �?                      �?              6@      �?      "@      �?                       @      @      �?      @      "@              ?@             �@@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ^�OQhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @���'@�	           ��@       	                   �4@"|z��@�           ��@                           �?MԮ���@E           ��@                            �?�i�o�@.           �~@������������������������       �ηP8�@�            �v@������������������������       �%
CG� @O             _@                            �?�`�ޗ<@            �@������������������������       �|~�ː@�            �q@������������������������       ��]��	@d           �@
                           @y��/�@�           T�@                          �<@运uÁ	@           �@������������������������       ��~dg[	@�           p�@������������������������       �����8�@c            �b@                          �6@� T�S@�           ��@������������������������       �b�V�{f@�            �n@������������������������       �y�P�ǁ@           �{@                           �?.�D�}�@�           ,�@                          �5@��JV�@�            @u@                           @%��1e+@|            �g@������������������������       ��G����@b            �b@������������������������       �(�"�>�?            �D@                           �?����S@V            �b@������������������������       ���j�6@:             [@������������������������       �]�$���?            �D@                          �9@W�:��@�           ��@                           @Y�\,b�@~           ��@������������������������       ���C�>n@$           `}@������������������������       ��>2�@Z            @_@                           �?*�m�q�	@r            �d@������������������������       ��n�ac�	@&             N@������������������������       �l���Y@L             Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     x�@      :@      G@      |@     @S@     ��@      m@     h�@     Pv@      ;@      $@     �i@     �x@      *@      8@     �r@     �L@     ��@      e@     �@      p@      4@             �P@      e@      @       @      ^@      "@     �~@     �P@     �q@     �Y@      @              5@     �R@              @      <@             �j@      3@     �X@      =@      @              2@      L@              @      8@             �a@      0@     �S@      8@       @              @      2@                      @             @Q@      @      4@      @       @             �F@     �W@      @      @      W@      "@     @q@     �G@      g@     �R@       @              *@      A@                     �C@      �?      W@      7@     �J@      <@       @              @@      N@      @      @     �J@       @      g@      8@     �`@      G@              $@     `a@     �l@      $@      0@      f@      H@     �p@     �Y@     pt@     `c@      ,@      $@     @Y@      [@       @      ,@     �Y@      B@     �X@     �R@      a@     �Y@      *@       @      T@     @X@       @      (@     @U@      7@      W@     �K@     �]@     �O@      (@       @      5@      &@               @      1@      *@      @      3@      2@     �C@      �?              C@     @^@       @       @     �R@      (@      e@      =@     �g@     �J@      �?              $@     �J@      �?      �?      <@      @      R@      @     �M@      (@                      <@      Q@      �?      �?      G@      @      X@      9@     ``@     �D@      �?      "@      V@     @d@      *@      6@     @c@      4@     @p@     �O@     @i@     �X@      @              9@      H@               @      F@             �\@      0@     �P@      2@                      "@      4@              @      *@             @V@      @     �D@      &@                      @      4@              �?      $@             �N@      @      B@      $@                       @                       @      @              <@              @      �?                      0@      <@              @      ?@              :@      &@      9@      @                      0@      ;@              @      8@              &@      &@       @      @                              �?                      @              .@              1@      �?              "@     �O@     �\@      *@      ,@     �[@      4@      b@     �G@      a@     @T@      @      @      C@      Y@      $@      *@     @X@      (@     �]@      ?@     �\@     �J@      @      @      A@     @U@      $@      *@     @U@      "@     @T@      >@     �S@     �B@      @              @      .@                      (@      @     �B@      �?      B@      0@      �?      @      9@      ,@      @      �?      *@       @      ;@      0@      5@      <@      @      @      "@      @              �?      @      @      @      @       @      (@      �?              0@      $@      @              @      @      7@      (@      *@      0@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$��ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��#׈S@�	           ��@       	                     �?�}�3i@           ֥@                           �?|�sn�@�           ��@                           �?�]X�.	@8           �|@������������������������       ���uF&�@~            @g@������������������������       �]�_H	@�            0q@                           @^z�W`V@y           �@������������������������       �11��8@z            @i@������������������������       ����c`�@�            0y@
                          �4@s�*WY�@P           �@                            �?>���@           0�@������������������������       �G�0�@G           (�@������������������������       �C��`@�            r@                           �?��=��@>           ،@������������������������       �K��L�U	@�            `q@������������������������       �tu�0#u@�           (�@                           �?ͳ~��@�           x�@                           �?���8)@@!           �{@                           @�?j��@m             e@������������������������       ��h(���@R            @^@������������������������       � L_^��?            �G@                           �?)[y��d@�            pq@������������������������       ����A��@e            @d@������������������������       �Y\�Xe@O            @]@                           �?�"	�9@�           ��@                          �3@O���@p            @e@������������������������       ���x�^ @3            �S@������������������������       �����@=            �V@                           @�#c�m	@9           P@������������������������       �
5<{C�	@G            �\@������������������������       ��j��@�             x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     �@      5@      M@     �}@     @T@     ��@      i@     �@     `w@      >@      *@     �k@     `x@      "@     �@@     �t@     �O@     H�@     �b@     Ё@     @o@      4@      @      Y@     �a@      @      "@     �^@      5@     �r@     �P@     @h@     @W@      ,@      @      L@     �Q@       @       @     �P@      .@      O@      F@     @S@      G@      (@       @      (@      :@              @     �B@       @     �B@      ,@      B@      (@      @      �?      F@      F@       @      @      =@      *@      9@      >@     �D@      A@       @              F@     @R@      �?      �?     �L@      @     @m@      7@     @]@     �G@       @              ,@      A@              �?      9@      @      L@      *@      C@      0@       @              >@     �C@      �?              @@      @     @f@      $@     �S@      ?@              $@     �^@     �n@      @      8@      j@      E@     |@     @T@     �w@     �c@      @      �?      G@     �Z@      @      @     �U@       @     �q@      >@     �e@     �O@       @      �?      @@     �Q@      @      @      L@      @     `d@      7@     �\@      E@      �?              ,@      B@                      >@      @     �]@      @     �M@      5@      �?      "@      S@     �a@      �?      3@     �^@      A@      e@     �I@     `i@     �W@      @       @     �@@     �F@      �?      &@     �C@       @      :@      <@      @@      G@      �?      �?     �E@      X@               @      U@      :@     �a@      7@     `e@      H@      @      (@     �V@     `c@      (@      9@     `b@      2@     �p@     �J@      i@      _@      $@      @     �@@     �K@       @      @      N@      @     @^@      "@     �U@      J@      @              *@      3@              @      0@             �P@      @      B@      &@                      *@      2@              @      &@             �C@      @      8@      $@                              �?              �?      @              ;@              (@      �?              @      4@      B@       @      @      F@      @     �K@      @      I@     �D@      @      @      0@      2@      @       @      B@      @      3@      @      5@      <@      �?              @      2@      �?      �?       @       @      B@       @      =@      *@      @      @      M@      Y@      @      2@     �U@      (@     �b@      F@     �\@      R@      @              .@      >@                      *@             �O@      &@      =@      "@                      @       @                       @             �C@      �?      3@      @                      "@      6@                      &@              8@      $@      $@      @              @     �E@     �Q@      @      2@     �R@      (@     �U@     �@@     �U@     �O@      @      @      (@      3@      �?      @      5@      @      $@      3@      &@      @      @      @      ?@     �I@      @      ,@     �J@      "@      S@      ,@     �R@      L@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��q9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�=$��/@�	           ��@       	                    �?���x@           ��@                           �?I���k�@6           P@                            @��o�@u            �g@������������������������       �@����@X            �a@������������������������       �Թ���*@             H@                            @\s�}@�            �s@������������������������       ���5p@8@b            @e@������������������������       �l'�^v�@_            �a@
                          �8@� �.S�@�           ȇ@                           @@�S�C� @�           @�@������������������������       �T˼�	@\             a@������������������������       ���H� @2           �@                          �:@��;���@J            @\@������������������������       ��(u��� @            �E@������������������������       ��oI���@/            �Q@                           @��[��@�           ��@                           @�Ȉ��@a           �@                           @��H�	@�           |�@������������������������       ��{(�@�           (�@������������������������       �kt���	@�           Ї@                           @�1#��@�           ��@������������������������       �s�����@�           �@������������������������       ���K�+@�            �p@                           !@�~['[	@0             S@                           �?�]�<P@"            �J@������������������������       ����ԹU@             5@������������������������       ��^Jϕ+@             @@                           @��D��@             7@������������������������       ��D=�U�@             (@������������������������       ��)���?             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     Pt@     ��@      ;@      K@      ~@     �Q@     ,�@      k@     �@     �s@      =@       @     �R@     `f@      @      $@     ``@       @     }@     �D@     �p@     �Q@      @       @      E@     �T@      @      @     @Q@              \@      =@     @Y@     �H@      @       @      (@     �@@                      ;@             �D@      @      I@      1@               @      &@      3@                      6@              >@      @     �B@      *@                      �?      ,@                      @              &@              *@      @                      >@     �H@      @      @      E@             �Q@      6@     �I@      @@      @              ,@      0@              @      :@              D@      *@      A@      1@      @              0@     �@@      @       @      0@              ?@      "@      1@      .@                      @@     @X@              @      O@       @     v@      (@     @e@      6@       @              @@     @U@              @      I@      �?     �s@      @     �`@      1@      �?              (@      2@              �?      4@             �H@       @      @@      @                      4@     �P@               @      >@      �?     �p@      @     �Y@      ,@      �?                      (@                      (@      @      A@      @     �A@      @      �?                      �?                      �?      @      ,@      �?      1@      @                              &@                      &@      �?      4@      @      2@       @      �?      2@     `o@     Px@      8@      F@     �u@      O@     Ё@      f@     0@     �n@      6@      ,@     �m@      x@      7@     �E@     �t@      L@     ��@     �d@     `~@     �n@      2@      *@      e@      n@      4@      :@     �n@      E@      i@     �`@     �l@     �d@      1@      "@     �S@     �Z@      @      1@     �`@      4@     �Z@      E@      ^@     �X@      @      @     �V@     �`@      ,@      "@     �[@      6@     �W@      W@     �[@     �P@      ,@      �?     @Q@      b@      @      1@     @V@      ,@     �v@     �@@      p@     �T@      �?      �?      J@      ]@              @      O@      @     0r@      .@     �g@     �N@      �?              1@      =@      @      $@      ;@      $@     �Q@      2@     @P@      5@              @      *@      @      �?      �?      ,@      @      @      "@      *@      �?      @      @      @       @      �?      �?      (@              @      "@      @      �?       @      @      @      �?                      @                       @       @      �?       @              @      �?      �?      �?      @              @      @      @                              @      �?                       @      @                      @               @               @      �?                      �?      @                      @               @              @                              �?      @                      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@O̼-:@�	           ��@       	                   �1@�T�@e           ̠@                           �?���;ڭ@�           ��@                           @L��3�@{            `i@������������������������       �TY�^@r             g@������������������������       �e>A:� @	             2@                           @7I. ���?           `z@������������������������       �P�=8��?�             j@������������������������       �ޤ�e� @�            �j@
                           �?9���Ȥ@�           ԗ@                           @$�%�@?           @������������������������       �J�Rx�@�            �r@������������������������       ��,V�?}            `h@                          �4@*��sׯ@�           �@������������������������       ���xD��@�           `�@������������������������       ������7@�             o@                            �?�1� l@f           ��@                           @�=	ݶ�@I           ��@                          �<@;���s	@r           ؁@������������������������       ��	�/vR	@"           @|@������������������������       �K��P�,@P            �]@                           @m��u
!@�            �u@������������������������       �?T6��R@�            �i@������������������������       ��=��@M            `a@                           @&t�V"�@           p�@                           @��<M�@�           ��@������������������������       ���u�@9           �}@������������������������       ����@�            �q@                          �;@�2��h@7            �U@������������������������       �xY8sL@,            �Q@������������������������       ���@             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     0s@     Ё@      >@     �H@     P{@      U@     Џ@     @h@     p�@     �x@      A@       @      ]@      t@      &@      9@      h@      B@     ��@      S@     �}@      e@      0@              7@      X@      �?      @      H@       @     �p@      ,@     �_@      D@      �?              .@      E@      �?              @@       @     �D@      @     �E@      5@                      (@      E@      �?              8@             �C@      @      D@      5@                      @                               @       @       @              @                               @      K@              @      0@             �l@       @      U@      3@      �?              @      ;@              �?      @             @`@      @      =@      @      �?              @      ;@               @      *@             �X@       @     �K@      *@               @     @W@      l@      $@      6@      b@      A@      {@      O@      v@      `@      .@              ;@     @P@      @      @      <@      @     `g@      &@     �`@      ?@                      8@      C@      @       @      8@      @     @S@      $@     �V@      :@                      @      ;@              @      @             �[@      �?      E@      @               @     �P@     �c@      @      1@      ]@      ;@     �n@     �I@     `k@     �X@      .@       @     �K@      \@      @      &@      T@      0@     �i@      E@     `c@     �S@      &@              &@     �G@      �?      @      B@      &@      D@      "@      P@      3@      @      @     �g@     @o@      3@      8@     �n@      H@     �s@     �]@     �r@     @l@      2@      @     @Z@     �^@      &@      *@     �_@      A@     `c@      P@     `a@     �`@       @      @      R@      T@      @      *@     �V@      =@      O@     �G@     �P@     @W@       @       @      O@      Q@      @      (@      T@      0@      M@      B@      I@      K@      @       @      $@      (@              �?      $@      *@      @      &@      0@     �C@      �?             �@@     �E@      @             �B@      @     @W@      1@     @R@     �D@                      5@      ;@      �?              1@      �?     �P@      *@      B@      8@                      (@      0@      @              4@      @      :@      @     �B@      1@              �?     �U@     �_@       @      &@     �]@      ,@      d@      K@     �d@      W@      $@      �?     �R@     @Z@       @      &@     �Y@      *@     �a@      H@     �c@      V@      @      �?     �Q@     �Q@      @      @     @T@      "@     �O@     �B@      P@      O@      @              @      A@      �?      @      6@      @      T@      &@     �W@      :@                      &@      6@                      .@      �?      2@      @      @      @      @              &@      3@                      $@      �?      .@      @      @       @      @                      @                      @              @              @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�N�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@Ly3�=@�	           ��@       	                    �?�Z���@�           N�@                           �?��w�@�           0�@                            @�c���@�            �k@������������������������       �>�wL�@N             _@������������������������       ���cJkS@C            �X@                            �?�����@R           8�@������������������������       ��uvv��@T            �a@������������������������       �5Ƨ2�@�            �y@
                          �1@�@�-@@�           ��@                          �0@�D�x?� @#           p|@������������������������       ��[$���?d             e@������������������������       �w�NO� @�            �q@                           @%�ЇV2@{           Ў@������������������������       ��O��@�           H�@������������������������       �i��{�@�            w@                           �?� t\(�@6           ��@                           �?��J�:�@"           �{@                           �?u��-��@�            @m@������������������������       ����_�@7            �V@������������������������       ��DX�H@_            �a@                           �?�y÷�m@�            @j@������������������������       ����q@G             ]@������������������������       �2���3@E            �W@                            �?N2HxU6	@           ��@                           @Ĳ�d"	@�           ��@������������������������       ��Nү�@N            �@������������������������       �������@A            �[@                           @/p�P0	@�           ��@������������������������       ��]���:	@           `{@������������������������       �u#�.��@y            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     �@      @@     �G@     `~@     �T@     \�@     @p@     8�@     �t@      4@      @     @\@     �s@      1@      6@     �m@      ?@     0�@     @Y@     �}@      c@       @      @      M@     �Z@       @      @     `a@      4@     `d@      L@      ^@     �T@       @              .@     �@@              �?      @@      �?     @R@      "@     �E@      .@      �?               @      2@                      7@             �A@      @      9@      "@      �?              @      .@              �?      "@      �?      C@      @      2@      @              @     �E@     �R@       @      @     �Z@      3@     �V@     �G@     @S@     �P@      @              *@      $@                      <@      "@      8@      (@      8@      0@      @      @      >@      P@       @      @     �S@      $@     �P@     �A@     �J@     �I@      @             �K@      j@      "@      .@     @X@      &@     �@     �F@      v@     �Q@                      *@     �P@              @      5@              l@      &@     �Y@      *@                      @      >@                      @             �U@              A@      "@                      $@     �B@              @      .@             @a@      &@      Q@      @                      E@     �a@      "@      &@      S@      &@     0v@      A@     @o@     �L@                      =@     �U@      �?      "@     �G@      @      n@      $@     �d@      7@                      *@      K@       @       @      =@      @     �\@      8@     �T@      A@              (@     `g@      m@      .@      9@     @o@     �I@     s@     �c@     �p@     `f@      (@      �?      E@     �J@      �?      @     �M@       @     ``@      9@     �X@      ;@      �?      �?     �A@      8@              @     �C@             �F@      3@     �F@      5@      �?      �?      2@      @                      *@              <@       @      2@      @      �?              1@      2@              @      :@              1@      1@      ;@      1@                      @      =@      �?              4@       @     �U@      @     �J@      @                      @      0@                      *@              J@      @      9@       @                      @      *@      �?              @       @      A@       @      <@      @              &@      b@     `f@      ,@      5@     �g@     �H@     �e@     �`@     �e@      c@      &@      @     @R@     �T@      @      ,@      W@      >@     �T@     �U@     �V@     @P@      @       @     @P@     @R@      �?      ,@     �S@      8@     @R@     �J@     @S@      J@      @      �?       @      "@       @              ,@      @      $@     �@@      *@      *@       @       @      R@     @X@      &@      @     �X@      3@     �V@      H@     �T@     �U@      @      @      P@      R@       @      @      P@      0@      F@     �C@     �F@     �Q@      @      �?       @      9@      @      @     �A@      @     �G@      "@      C@      1@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�J/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @'e�n4@�	           ��@       	                    �?�(|Sb�@�           j�@                            �?pI��@           ��@                          �5@H���o@=            �@������������������������       �A⭕�@�            �o@������������������������       �<���ɮ	@�             p@                          �;@ƵD_�@�           ��@������������������������       �]�K6�@^           ��@������������������������       �ъD��@�            �g@
                            @���V�@u           �@                            �?l���	�@           0y@������������������������       ��$���@�            Ps@������������������������       ��6 ~��@:            �W@                           �?�;n��@n            @e@������������������������       ���uGV@            �F@������������������������       �I�o+d�@S            @_@                           @C�`�(E@8           P�@                           @L*B��@�           �@                            @��o�W@�           ��@������������������������       �D��or�@U           ��@������������������������       �=#Gv��?\            �b@                          �<@:e?�x@.            }@������������������������       ��84�k@            {@������������������������       �ǒY��_@             @@                          �4@2q>���@Y             c@                          �1@�D� �c@#            �L@������������������������       ���l����?             &@������������������������       ��ПK)@             G@                          �6@Ж�h�@6            �W@������������������������       �v��d�@             9@������������������������       �ڤhne@(            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     x�@     �@@      L@     �}@     �Q@     $�@     �h@     ��@     �t@      B@      1@     �k@     �u@      5@     �@@     �s@      M@     �w@     �d@     @z@     �k@      :@      1@     �d@     �p@      3@      :@     �o@     �G@     �n@     �]@     �r@     @f@      8@      @     �F@     @S@      @      "@     @T@      *@     @V@      G@     �X@      C@      "@              4@     �C@                     �A@      �?      L@      6@     �N@      .@      @      @      9@      C@      @      "@      G@      (@     �@@      8@      C@      7@      @      ,@      ^@     �g@      0@      1@     �e@      A@     `c@     @R@     �h@     �a@      .@      @     @X@     �d@      *@      *@     �b@      9@      b@      O@      f@     �V@      ,@       @      7@      8@      @      @      5@      "@      &@      &@      7@      I@      �?              M@     �S@       @      @      P@      &@     @a@     �F@     �^@     �F@       @             �B@     �G@              @     �H@      $@      X@     �@@     @X@      ;@       @              =@      G@              @      @@       @      Q@      6@      T@      1@       @               @      �?                      1@       @      <@      &@      1@      $@                      5@      @@       @       @      .@      �?      E@      (@      9@      2@                      @       @                      "@              .@      �?      *@       @                      2@      >@       @       @      @      �?      ;@      &@      (@      0@              �?     �S@     �j@      (@      7@      d@      *@     X�@     �A@     �w@     @[@      $@      �?      P@     @g@      @      4@     �a@      "@     x�@      ?@      v@     @W@      @      �?     �D@     @b@              @     �W@      @     P|@      &@     `o@     �M@      �?      �?      >@     �`@              @     �T@      @      x@      &@     `i@     �M@      �?              &@      (@                      &@      �?     �P@              H@                              7@      D@      @      *@     �H@      @     @e@      4@     @Y@      A@       @              7@      D@      @      *@     �C@      @      e@      1@     @W@      9@       @                                              $@      �?      �?      @       @      "@                      .@      <@      @      @      2@      @      <@      @      8@      0@      @              �?      &@              @       @              *@              ,@      *@                                              @                      @               @       @                      �?      &@                       @              "@              (@      &@                      ,@      1@      @              0@      @      .@      @      $@      @      @                              @              @       @      @               @              @              ,@      1@                      (@       @      "@      @       @      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�S-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���W߀@�	           ��@       	                   �4@ϊ���@�           ��@                           �?)Pz��N@8           H�@                           �?�Wt�s�@�            `s@������������������������       �"�L81@R            @a@������������������������       ��WKH��@j            �e@                          �1@\���2@|           ��@������������������������       �}-B�S�@n            @e@������������������������       ���nN/g@           �z@
                            @���	@H           D�@                           �?���	@�           X�@������������������������       ���C1K*	@�            �s@������������������������       ��:�8�	@2           0@                          �?@b4���1	@Q           0�@������������������������       ��G�q��@;           �@������������������������       �D���@            �C@                           @x77S��@           ��@                           �?xT�@�           ��@                          �4@Bj��?�            pv@������������������������       �jĀ��b�?�             m@������������������������       ���Y�@O            �_@                            �?����.�@�           �@������������������������       �ο6��D@m             e@������������������������       ��0n��@           Ђ@                          �7@����Z�@E           0�@                           @��x9�@�            �u@������������������������       �>���8@�            0q@������������������������       �y�q�@&            �Q@                           �?��;o@k            �e@������������������������       �D�GrW�?"             K@������������������������       ����O@I            �]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@      s@     �@      <@      O@     �~@     �T@      �@     �i@     ��@     �u@     �C@      5@      m@     �v@      3@      H@     pu@     �P@     @v@      e@     @w@     `n@      B@      @     �N@     @`@       @      ,@     �a@      &@     �i@     �P@     �g@     �Q@      @              0@      G@              @      B@      �?     �U@      ,@     �V@      ,@      �?              @      ,@               @      9@      �?      A@      *@      C@      @      �?              (@      @@              @      &@             �J@      �?      J@       @              @     �F@      U@       @      "@      Z@      $@     @]@      J@     @Y@      L@      @              .@      @@       @      �?      ,@      @      E@      ,@      @@      .@              @      >@      J@      @       @     �V@      @     �R@      C@     @Q@     �D@      @      1@     �e@     �l@      &@      A@     `i@     �K@      c@     �Y@     �f@     �e@      >@       @     �Y@     �\@      @      :@      ^@     �@@     �U@     @Q@      ^@      [@      2@      �?      E@     �I@      @      @     �F@      .@     �@@      =@      ?@     �I@      @      @     �N@     �O@       @      5@     �R@      2@      K@      D@     @V@     �L@      (@      "@     @Q@     @]@      @       @     �T@      6@     @P@     �@@     �N@     @P@      (@      @     @P@     �[@      @      @     @S@      6@     @P@      >@      K@      O@      (@      @      @      @       @      @      @                      @      @      @                     �Q@      k@      "@      ,@     �b@      0@      �@     �C@     �y@     @Z@      @             �H@     `b@       @      @     �V@      &@     �|@      8@     pq@      O@      �?              &@     �H@                      3@      @     �h@      @     �Q@      @                      @      <@                      @             `b@      �?     �G@                              @      5@                      ,@      @     �H@      @      8@      @                      C@     �X@       @      @      R@       @     �p@      3@      j@     �L@      �?              .@      5@       @              (@             �Q@       @      =@      1@                      7@     @S@              @      N@       @     @h@      1@     `f@      D@      �?              6@     �Q@      @      &@     �M@      @     �b@      .@      a@     �E@       @              (@      L@      @      @     �D@      @     @^@      @     @S@      3@       @              $@      E@              @      ?@      @     �Y@      @     @Q@      &@      �?               @      ,@      @      @      $@              3@               @       @      �?              $@      ,@       @      @      2@       @      ;@      (@     �M@      8@                              @                      @              0@              9@      @                      $@       @       @      @      .@       @      &@      (@      A@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��./{@�	           ��@       	                     @c�e��@           �@                           �?不���@*           ��@                           �?��x+�@�            `r@������������������������       �$�h�W@N            �]@������������������������       ��1����@k            �e@                           �?ʯ��@q           ȁ@������������������������       �5�9.� @�            �s@������������������������       �6��eM@�            �o@
                           @�$��@�            pv@                           �?;� �l�@�            p@������������������������       ��Z��k@"             I@������������������������       ��˚M�@y            �i@                           @X�����?>            �Y@������������������������       �RA"]�?             <@������������������������       �n`�*V�?-            �R@                          �3@>vRhS@�           �@                           @�Y�@A           Ȍ@                          �1@D2b�%�@}            �@������������������������       �`=D�IC@�            `p@������������������������       �:ЏQ!@�            �u@                          �0@�$���@�            �s@������������������������       ����2! @            �J@������������������������       �RlrO�@�            @p@                            �?�S.� 	@`           ��@                           �?�h�5�@4           �~@������������������������       ��T���@             i@������������������������       ��މ	@�            Pr@                          �9@YV,�'	@,           ��@������������������������       ��W��x@-           `�@������������������������       �T+�0�	@�            y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     x�@     �C@      M@     �}@     �S@     P�@      l@     Ї@     �w@      ?@              R@     �d@      @      (@     �^@      $@     �{@      @@     `o@     @X@      "@             �H@      `@       @      @     @T@      $@     Pt@      6@     �e@      M@      "@              5@     �E@       @      @     �G@             @Q@      (@      L@     �A@      @              $@      &@       @      @      3@              <@       @      1@      4@      �?              &@      @@              �?      <@             �D@      @     �C@      .@      @              <@     @U@               @      A@      $@      p@      $@     @]@      7@      @              *@     �E@               @      4@      @     @d@      @      N@      "@                      .@      E@                      ,@      @     �W@      @     �L@      ,@      @              7@      B@      @      @     �D@             �^@      $@     �S@     �C@                      4@      A@      @      @     �B@              O@      "@      G@     �C@                      @      @                       @              :@      �?      @      @                      .@      <@      @      @     �A@              B@       @     �C@      B@                      @       @                      @              N@      �?      @@                              �?      �?                                      $@              0@                               @      �?                      @              I@      �?      0@                      5@      j@     �x@     �@@      G@     @v@      Q@     X�@      h@     �@     �q@      6@      @      J@     �`@      @      @      X@      @     �p@     �I@     `i@     @V@      @      @      ?@      S@      @      @      R@      @      e@     �@@     �b@     �N@                       @      <@               @      6@              U@      "@     �T@      ;@              @      7@      H@      @      @      I@      @      U@      8@      Q@      A@               @      5@      L@       @       @      8@      �?     �Y@      2@     �J@      <@      @              @      $@                      �?              ;@              @      @               @      1@      G@       @       @      7@      �?     �R@      2@     �G@      7@      @      0@     �c@     pp@      <@     �C@     @p@     �N@     �q@     �a@     @s@     @h@      2@              M@     �Q@      @      $@      S@      0@     �R@     �N@     �R@      G@      @              :@     �D@      �?              A@      �?      7@      =@      =@      .@      �?              @@      =@       @      $@      E@      .@      J@      @@     �F@      ?@      @      0@     �X@      h@      9@      =@      g@     �F@     @j@     @T@     @m@     �b@      ,@      @      O@     �a@      ,@      3@     �`@      :@     �d@     �G@     �e@     �R@      ,@      &@      B@      J@      &@      $@     �H@      3@      F@      A@     �N@     �R@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ+�]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �1@G��ˇX@�	           ��@       	                    �?{ d@�@�           X�@                           �?'<��+�@z            `h@                            �?4~�mR@5            �T@������������������������       ���=�@             B@������������������������       �K7i�P�@             G@                           �?�΁� @E            @\@������������������������       ��1���@            �E@������������������������       ��l��8�@+            �Q@
                           @lۧ�3 @           �|@                            �?%��|�|�?�             w@������������������������       �������?8            @X@������������������������       �F�u� @�            �p@                          �0@ťY�r�@5             V@������������������������       � ��] @             =@������������������������       ����yT @%            �M@                            �?��)��@           |�@                           @����&�@)           X�@                           �?K��f1�@h           ��@������������������������       ����xW@�            �i@������������������������       ��x#9D�@�            `v@                           @t߹L!�@�            �s@������������������������       �$�'�<h@1             S@������������������������       ���m�@�            �m@                            @����@�           ��@                            �?l^��A�@}           |�@������������������������       ��0�	�G@           ��@������������������������       �㶸�8@b           @�@                           �?ܮ��E|@_           ��@������������������������       ��c)�i@�            Pq@������������������������       ��M^�$X	@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     ps@     p�@      @@     �I@     `{@      X@     �@     @j@     ؈@     u@      @@              <@     �X@      �?      @      C@       @     �p@      7@     �b@      C@      �?              .@     �B@      �?       @      8@       @     �D@      (@     �C@      6@                      @      $@      �?              &@       @      6@      @       @      1@                      �?      "@                       @       @      @      @      @      "@                      @      �?      �?              "@              1@      @      @       @                      &@      ;@               @      *@              3@      @      ?@      @                              @                      @              "@      @      2@      @                      &@      5@               @      "@              $@       @      *@       @                      *@     �N@              �?      ,@             `l@      &@      \@      0@      �?              *@      I@                      @              h@      @     @V@      $@                              "@                                     �P@      @      0@      @                      *@     �D@                      @             �_@      @     @R@      @                              &@              �?      @             �A@      @      7@      @      �?                       @                       @              &@               @      @                              @              �?      @              8@      @      5@              �?      6@     �q@     �|@      ?@      H@      y@     �W@     ؇@     `g@      �@     �r@      ?@       @      U@      ]@      @      *@     @X@     �@@     @k@     �P@     �e@     �N@       @       @     �O@     @S@       @      *@     �Q@      :@     @X@      K@     �[@      D@       @              7@     �@@      �?       @     �@@      $@      D@      5@      :@      (@      @       @      D@      F@      �?      &@     �B@      0@     �L@     �@@     @U@      <@      @              5@     �C@      @              ;@      @     @^@      (@     �N@      5@                      &@      (@       @               @              =@      @       @      @                      $@      ;@      �?              9@      @      W@      @     �J@      .@              4@     �h@     �u@      :@     �A@     �r@     �N@     �@     @^@     �}@     �m@      7@       @     @\@      i@      .@      ,@      g@     �C@     �u@      R@     0r@     @a@      *@      @      R@     �_@      *@      $@     �W@      <@     �g@      G@     �d@     @W@      &@       @     �D@     �R@       @      @     @V@      &@     `d@      :@      _@     �F@       @      (@     �U@     �a@      &@      5@     �]@      6@     @h@     �H@     �f@      Y@      $@              7@     �E@              @      2@              W@      &@     �P@      0@              (@     �O@      Y@      &@      ,@     @Y@      6@     �Y@      C@     �\@      U@      $@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�PpyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Ωs� E@�	           ��@       	                   �6@G��\�@           ��@                            �?ۥ��0@!           0�@                           @�X��K~ @�            �l@������������������������       ��`
rL@F            �^@������������������������       �4OM	���?B            �Z@                            �?��H��@�           �@������������������������       �3����u@�            @n@������������������������       ��S�#G@�             y@
                            @���*�@�            �w@                            �?A�@�            �p@������������������������       �����D@�            @i@������������������������       ����z�a@*            �O@                           @*�W/&~@C            @\@������������������������       ��ҦSt@7            �W@������������������������       �Њ���r�?             3@                           �?Q��� @�           Ҥ@                           @����	@~            �i@                          �8@�c�	�@T            `a@������������������������       ��)�
@6             V@������������������������       �������@            �I@                            @�G��@*            �P@������������������������       ���!�p@#             J@������������������������       ��\�>��@             .@                           @%��@           6�@                          �6@���ޢ@�           ��@������������������������       �����3@�           �@������������������������       ��z���@J           x�@                           !@��<��j	@4            �T@������������������������       ������@%            �M@������������������������       �c���@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `r@     ��@      @@     �L@     �z@     �Q@     ,�@     `m@     (�@     pw@     �@@      @     @S@     �c@      @      *@     �[@      @     @{@     �J@     �r@     �T@       @             �H@     �Z@               @      N@      @     0v@      :@      j@     �J@       @              @      7@              �?      &@             �Y@      @     �Q@      *@                      @      ,@              �?      &@              >@      @      J@      @                              "@                                      R@              2@      @                     �F@     �T@              @     �H@      @     �o@      6@     @a@      D@       @              2@     �E@              @      3@             �S@      "@      M@      (@       @              ;@      D@              @      >@      @     �e@      *@      T@      <@              @      <@      I@      @      @     �I@      @     @T@      ;@     �V@      >@      @      @      7@      D@       @      @      =@      @     �I@      *@     �P@      9@      @      @      0@      ;@       @      @      9@       @     �B@      *@     �H@      3@      @              @      *@                      @       @      ,@              1@      @                      @      $@      �?       @      6@              >@      ,@      8@      @                      @      $@      �?       @      6@              1@      &@      5@      @                                                                      *@      @      @                      .@      k@     pw@      =@      F@     �s@     �O@     ��@     �f@     �@     @r@      9@      @      6@      9@              @     �D@       @      5@      ;@      =@      3@              @      5@      ,@              @      =@      @      @      4@      .@      0@              @      "@      "@              @      8@       @      @      @      *@      (@              @      (@      @              @      @       @              ,@       @      @                      �?      &@                      (@      @      .@      @      ,@      @                      �?      $@                      $@       @      *@       @      (@       @                              �?                       @       @       @      @       @      �?               @     `h@     �u@      =@     �B@     @q@     �K@     �@     `c@     �}@     q@      9@      @     @g@     �u@      ;@     �A@     `p@      H@     ؁@     �`@     `}@     �p@      8@       @     �W@     @j@       @      ;@      a@      4@     �{@      Q@     �s@     �`@      @      @      W@     �`@      3@       @     @_@      <@      `@     �P@     �b@      a@      1@       @      "@      @       @       @      ,@      @      @      4@       @      @      �?       @       @      @       @       @      $@              @      1@      @      @                      �?       @                      @      @              @      @       @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJW`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�^�@�	           ��@       	                    @�)�^��@{           ��@                           �?Nh� �6@E           ��@                           �?M���s@�            �s@������������������������       �Q�EҴ@=            @Y@������������������������       ��T�;L@�            �j@                           �?Y�#�@�           �@������������������������       �;67��J@�            py@������������������������       �vu���@�            �i@
                          �1@
���۪ @6           8�@                          �0@&1���?�            0v@������������������������       ��닳���?J             ^@������������������������       ���-���?�            `m@                           @i���@_            �@������������������������       �&�0�@M            @\@������������������������       �����7@           0{@                           �?[݈���@7           H�@                           �?R-���@u           �@                            �?�/�T�@�            @s@������������������������       ���龢'@j            `e@������������������������       �O�����@X             a@                          �=@Z�� m�@�            �p@������������������������       ����-@�            `n@������������������������       ����{4@             <@                           @u��!	@�           ��@                           �?s�i��	@U           X�@������������������������       �Uc�@k@>            �X@������������������������       ���*(�	@           @�@                           @+���@m           ��@������������������������       �9�4��@_           �@������������������������       ���}��9@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �p@     P�@      ;@     �H@      }@     @R@     ��@     �k@     ��@     @t@      B@      @      U@     �o@      @      .@     �d@      .@     H�@      T@     �z@     �]@      "@      @      K@     �a@      @      $@     @`@      &@     �j@      Q@     �g@      U@      "@              6@      C@               @      A@      @     @Z@      @     �S@      8@      �?              @      .@                      &@             �A@      �?      @@      @                      3@      7@               @      7@      @     �Q@      @     �G@      4@      �?      @      @@     @Z@      @       @      X@      @     �[@      O@      \@      N@       @      @      <@     �L@      @      @      S@      @     �L@     �A@     @T@     �G@       @              @      H@       @      @      4@      �?     �J@      ;@      ?@      *@                      >@      \@      �?      @      B@      @      {@      (@     `m@      A@                      @      E@              �?      *@             �h@      @     @U@       @                              4@                      @              Q@              5@      @                      @      6@              �?      "@             @`@      @      P@      �?                      9@     �Q@      �?      @      7@      @     �m@      "@     �b@      :@                      $@      ;@                      @      @      C@      @      ;@       @                      .@     �E@      �?      @      4@      �?     �h@      @     �^@      8@              0@     �f@     �t@      4@      A@     �r@      M@     �v@     �a@     @y@     �i@      ;@              H@     �\@      @      @     �O@      �?      b@      <@     @`@     �B@      @              >@      J@      @      @      @@      �?     �S@      &@     �R@      6@                      7@      7@      @              1@      �?     �D@       @      C@      1@                      @      =@              @      .@              C@      @     �B@      @                      2@     �O@               @      ?@             @P@      1@     �K@      .@      @              1@      O@                      :@              O@       @      K@      *@      �?              �?      �?               @      @              @      "@      �?       @      @      0@     �`@      k@      1@      =@     �m@     �L@     �k@     @\@      q@      e@      6@      0@     �X@     `b@      .@      4@     �c@     �G@     �U@     �V@     @^@      ^@      4@      @      ,@      (@              @      <@       @      @      ,@      @      @      @      $@     @U@     �`@      .@      .@     @`@     �F@     @T@      S@     �\@     @]@      1@              A@     @Q@       @      "@     �S@      $@      a@      7@      c@     �H@       @              <@     @Q@      �?      "@      S@      @     �`@      5@      c@     �H@       @              @              �?              @      @       @       @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����@�	           ��@       	                   �:@x+r1��@z           ^�@                           �?\�ojv@|           |�@                            �?i�U>�P@�           ȅ@������������������������       �h)�/@�            `k@������������������������       �6�6�o@3           �}@                          �8@��"�&T@�           ��@������������������������       �ע��$@o           0�@������������������������       �Vul��E@T             `@
                          �?@�����	@�             y@                            �?��;��k	@�            t@������������������������       ��&Ozy�	@7            �W@������������������������       �؈��@�            @l@                           �?��v-Z+	@1            �S@������������������������       ������b@             4@������������������������       �x�~��@%            �M@                          �7@
�g`j@2           h�@                           �?Hm�CS@9           ē@                           @ �A{z @           0{@������������������������       ������?�            �r@������������������������       ��!�l��@Z            �`@                           �?�2g�z@           ��@������������������������       �E|{�@           py@������������������������       �ɍ��h�@
           pz@                          �<@V=_p@Q@�            �z@                          �8@J���@�            �t@������������������������       �{e&�l@>             [@������������������������       �J�@PO@�            `l@                           @7��=
@6            �V@������������������������       �A��9��@             @@������������������������       �cx�x�@"             M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     0s@     P�@      =@      K@     �~@     �R@     ��@     �l@     ��@     `v@      C@      9@     �i@     �t@      7@      C@     �u@     �K@     0w@     �g@     �v@     �n@      ?@      @      e@     �q@      3@      <@     �q@      E@     �t@     �b@     �s@     �e@      :@              P@     �\@      (@      @      ]@      1@      a@     �P@     @T@      R@      $@              4@      :@      �?      @     �D@      @     @P@      3@      2@      1@      @              F@     @V@      &@      @     �R@      ,@      R@      H@     �O@     �K@      @      @     @Z@     �d@      @      6@     @e@      9@     @h@     �T@      m@      Y@      0@      @      X@     �a@      @      3@     �b@      9@     �e@     @P@     �j@     �W@      @              "@      8@       @      @      3@              5@      1@      2@      @      $@      2@      C@     �I@      @      $@      N@      *@      D@      D@      H@     @R@      @      *@      :@      E@       @      @     �G@      $@      D@      >@      F@      M@      @       @      @      *@       @       @      1@      @      $@      &@      1@      "@       @      &@      5@      =@              @      >@      @      >@      3@      ;@     �H@       @      @      (@      "@       @      @      *@      @              $@      @      .@      �?              @      @              @      @                      �?       @                      @       @      @       @               @      @              "@       @      .@      �?              Y@     �k@      @      0@      b@      4@     X�@     �C@      {@     @\@      @             @P@     �e@      @      $@     �U@      0@     �@      .@     @s@      S@      @              0@      K@      �?       @      7@      �?     �k@      @     @X@      *@      �?              (@     �A@                      .@      �?      e@             �N@      @                      @      3@      �?       @       @              K@      @      B@      @      �?             �H@     �]@      @       @      P@      .@     �q@      &@     `j@     �O@      @              ;@      O@       @      @     �E@      @      `@       @     �W@      ?@      �?              6@     �L@       @      @      5@      &@     @c@      @      ]@      @@       @             �A@      I@      �?      @      M@      @     @T@      8@     �_@     �B@      @              7@     �@@      �?      @     �E@      @     �P@      8@      [@      8@      @              ,@      $@                      1@       @      8@       @      ;@      "@      @              "@      7@      �?      @      :@       @     �E@      6@     @T@      .@                      (@      1@              �?      .@              ,@              2@      *@                      @       @              �?       @              @              $@      @                      @      .@                      *@              @               @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Y��c@�	           ��@       	                   �;@�:����@z           ��@                           �?C��p�\@�           @�@                          �3@ 4�=J@l           ��@������������������������       �����@�            p@������������������������       �gGA(4@�            `u@                           �?�iɉ	@L           �@������������������������       ���u�qQ	@^           (�@������������������������       �=����@�            @w@
                           @�%>M��	@�            s@                           �?'.y�p�	@�            �p@������������������������       �e�t	ޞ	@�             m@������������������������       ��Ō�3@            �B@                          �=@`�+��@            �A@������������������������       �7�FikN@
             2@������������������������       �	�O�@	             1@                           @c��<@/            �@                           @x�'\ϻ@�           $�@                           �?���8�@           pz@������������������������       ��T�	�) @T             `@������������������������       ���KK��@�            `r@                          �4@�?�_�@�           �@������������������������       ����Ԁ @#           �{@������������������������       �7����@�            `r@                           @԰}$��@H           �@                            @�}��>@1           �}@������������������������       �~}�V�T@�            Pv@������������������������       ���8R�N@H             ]@                           �?�pO��@             C@������������������������       �PK��@
             3@������������������������       ���\p�2@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �q@     ��@      B@      N@     p~@      V@     \�@     �m@     h�@     �u@      <@      *@     `i@     �s@      9@      F@     @v@     �O@     `z@     �h@     �t@     @o@      8@       @      f@      q@      2@      >@     pr@      H@     @y@     `e@     �r@      h@      4@              I@     �S@       @      @      Q@       @      i@      ,@      _@      G@       @              1@      @@                      :@      @     @U@      $@      K@      =@                     �@@      G@       @      @      E@      @     �\@      @     �Q@      1@       @       @     �_@     �h@      0@      7@     `l@      D@     �i@     �c@     �e@     @b@      2@       @     @X@     �`@      ,@      0@     �f@     �@@     �_@     �[@     �_@     @Y@      2@              >@      P@       @      @      F@      @     �S@     �G@      H@     �F@              @      :@      C@      @      ,@     �N@      .@      2@      ;@      @@      M@      @      @      :@      ?@      @      ,@     �J@      &@      .@      6@      >@      K@      @      @      4@      :@      @      ,@     �C@      $@      (@      3@      ;@     �J@      @              @      @                      ,@      �?      @      @      @      �?      �?       @              @                       @      @      @      @       @      @              �?              @                      @              @       @       @       @              �?              @                      @      @              @               @                     �T@     @o@      &@      0@     ``@      9@     ��@     �D@      x@      Y@      @              M@      d@       @      @     �T@      *@     �~@      3@     �p@      N@       @              <@      S@                      ;@      *@     �c@       @     �W@      3@      �?              @      :@                       @      �?      N@       @      >@      @                      8@      I@                      9@      (@      X@      @     @P@      .@      �?              >@      U@       @      @      L@             �t@      &@      f@     �D@      �?              ,@      H@       @       @      8@             `m@      @     @X@      3@                      0@      B@              �?      @@             �X@       @     �S@      6@      �?              9@     �V@      "@      *@      H@      (@     �`@      6@     �\@      D@       @              5@     �U@      @      (@     �D@      &@     �`@      *@      [@      D@       @              3@      S@      @      "@      @@      $@     @U@      "@      V@      6@       @               @      $@       @      @      "@      �?     �G@      @      4@      2@                      @      @       @      �?      @      �?      @      "@      @                              �?                      �?      @              @      @       @                              @      @       @               @      �?               @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJX�g7hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Ts�|X@�	           ��@       	                    �?ǿ4S�@x           ��@                          �;@�04-@�           ��@                           �?G����@�           H�@������������������������       ����L�>@�            q@������������������������       ��D$g�c@�            �u@                            �??�"`��@6            �S@������������������������       �����@             0@������������������������       ���~���@+             O@
                           �?h���Ce	@�           h�@                          �2@�g�r��	@�           �@������������������������       ��H��@~            �j@������������������������       ����F
@F           `�@                          �5@�V�t�@�            �y@������������������������       ���	KsZ@�            �l@������������������������       ���/���@l            @f@                           @���'@2           ��@                           @F�pu�@�           T�@                           �?�d޽PK@!           ȉ@������������������������       �C���D@�             t@������������������������       ��8�X�@K           p@                           �?`{�3� @�            �q@������������������������       ��V`�[��?.            @Q@������������������������       �.P���@�            �j@                          �3@�M(�(@Y           �@                           @+��U�T@�            `j@������������������������       ��fJ��^@e            �d@������������������������       �E3AŝB@             F@                          �7@�p�a�*@�             u@������������������������       �2I/��@n            �d@������������������������       �*-%���@j             e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     ps@     0�@      A@     �K@     �}@     �Q@     @�@     �k@     ��@     �v@      ;@      3@      l@     pu@      :@     �B@     pt@      H@     �w@     �g@      x@     p@      8@             �Q@     @Z@      @      @     @V@      @      e@     �B@     �b@      O@                      N@      W@      @       @     �Q@       @      d@      ;@      b@      K@                      ?@      @@      @       @     �F@      �?     @S@      .@      F@      6@                      =@      N@                      :@      �?      U@      (@      Y@      @@                      $@      *@              @      2@       @      @      $@      @       @                      @      @                      @       @                      @      �?                      @      $@              @      .@              @      $@      @      @              3@     `c@     �m@      6@      @@     �m@      F@      j@     �b@     `m@     `h@      8@      3@     �^@     �c@      2@      ;@     �f@      B@     �`@      _@      d@     �c@      5@      @      0@      5@              �?      G@       @      A@      :@      G@      2@              .@     �Z@      a@      2@      :@     �`@      A@     �X@     �X@     �\@     `a@      5@             �@@     @T@      @      @      M@       @     @S@      ;@     �R@      C@      @              @     �G@      @      @      =@      @      K@      .@      G@      7@                      <@      A@               @      =@      @      7@      (@      <@      .@      @       @     �U@     �i@       @      2@      c@      7@     x�@      @@     �x@     �Y@      @       @     �J@     �a@      @      @      X@      (@     �|@      *@     �p@      M@      �?       @      I@     �W@      @      �?     �R@      (@     `u@      *@     �g@      F@      �?       @      2@      F@                      .@       @     �d@      @     �K@      "@                      @@     �I@      @      �?     �M@      @     �e@      "@     �`@     �A@      �?              @     �F@              @      6@             �\@             �T@      ,@                              "@                      @             �D@              ,@      �?                      @      B@              @      2@             @R@             @Q@      *@                     �@@     �P@      @      ,@      L@      &@     �d@      3@      `@     �F@       @              .@      &@              @      8@             �S@      @     �L@      .@                      $@      &@              @      .@             �P@      @     �I@      @                      @                       @      "@              *@              @      "@                      2@      L@      @       @      @@      &@      V@      .@     �Q@      >@       @              @      C@      @      @      ,@      @     �H@              >@      *@       @              *@      2@              @      2@      @     �C@      .@     �D@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Zc%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�vO�/X@�	           ��@       	                     �?N�ӄ��@V           ��@                          �5@=��ӹ@�           P�@                          �1@h*�g#@�             s@������������������������       ��@�t�@,            @R@������������������������       �o�=�?!@�             m@                          �8@��� 
@�            �u@������������������������       �[f����@a             d@������������������������       �1R���
@s            �f@
                           �?o�S���@�           ė@                          �1@�{�&	@�           p�@������������������������       ��A�W�,@O            �^@������������������������       ��Dbu|r	@w           �@                          �3@�̱��@�            Py@������������������������       �٬l?��@\             a@������������������������       �/#�'iR@�            �p@                           �?�zl�@4           8�@                          �4@�֞���@i           0�@                          �0@M[m���?�             v@������������������������       �6�����?!             L@������������������������       �|������?�            �r@                           @k��ڗ@�            �l@������������������������       �<�d�?�@#            �O@������������������������       �es�x�@n            �d@                           �?���@�            �@                            @�ޭ�@_           Ё@������������������������       ��pԇ�i@+           �}@������������������������       �X�;@4             W@                           @�K��(@l           p�@������������������������       �3�� u@L            �a@������������������������       ��dC���@            |@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     �@      9@     �H@     �@     �W@     ��@      l@     �@     �u@      >@      1@      k@     �r@      3@      C@     `x@     �O@      w@     �f@     �s@     �m@      ;@      @     �Q@     �R@       @      *@      _@      3@     @^@     �L@     �V@     �M@      .@              7@      >@              �?     �P@      @     �R@      5@      M@      :@      �?              @      @                      @      �?      =@      @      0@       @                      1@      8@              �?     �O@      @     �F@      2@      E@      2@      �?      @      H@      F@       @      (@     �L@      ,@     �G@      B@     �@@     �@@      ,@              ;@      1@      �?      $@      >@      �?      =@      $@      2@      (@      @      @      5@      ;@      �?       @      ;@      *@      2@      :@      .@      5@       @      *@     @b@      l@      1@      9@     �p@      F@      o@     @_@     �k@     @f@      (@      *@     @Z@     @e@      0@      6@     @j@     �C@     �d@      V@      b@     �`@      (@      �?      @      5@                      <@              C@      @      0@      $@              (@     �Y@     �b@      0@      6@     �f@     �C@     �_@     �T@      `@     �^@      (@             �D@     �K@      �?      @      L@      @     @U@     �B@     @S@     �F@                      "@      3@                       @              C@      1@      =@      0@                      @@      B@      �?      @      H@      @     �G@      4@      H@      =@               @     �X@     �j@      @      &@     �^@      ?@     h�@      E@     P|@      [@      @              4@     �U@      �?       @      =@      &@     �p@      @     �a@      4@       @              &@      E@               @      (@             �g@       @     �T@      $@       @                      1@                      @              4@              *@      @                      &@      9@               @      "@              e@       @     �Q@      @       @              "@     �F@      �?              1@      &@     �S@       @     �L@      $@                       @      ,@                      (@       @      4@              @                              @      ?@      �?              @      @      M@       @      I@      $@               @     �S@     @_@      @      "@     �W@      4@     0x@      C@     �s@      V@      �?       @     �D@     �O@      @      @      P@      @     �f@      (@      b@     �G@      �?       @      C@      L@       @      @      L@      @     �b@      (@      \@      C@      �?              @      @      �?      �?       @              ?@              @@      "@                     �B@      O@       @       @      >@      0@     �i@      :@      e@     �D@                      "@      .@      �?      �?      @      &@     �E@      .@      =@      $@                      <@     �G@      �?      �?      7@      @     @d@      &@     �a@      ?@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Y�.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����@z	           ��@       	                    �?.��h-�@^           �@                          �;@42�/�@�           �@                           �?�Xo��Z@;           ��@������������������������       �;�l��J@           @z@������������������������       ���9/�@8            �@                            @5���v	@�            pq@������������������������       ��ͨݙ@a            `b@������������������������       ����g	@H            �`@
                           �?��
Q+@z           p�@                          �6@rÁ�6@�            �n@������������������������       �>P�\�9@a             b@������������������������       �Z<�@=            �Y@                            �?殏�?�@�            pu@������������������������       ���d�O@E            �Y@������������������������       �_��nV�@�             n@                           �?��?��@            �@                            �?r����M@d            �@                           �?NL��v�?Q            �a@������������������������       ��P�,�r�?&            @P@������������������������       �5��,�?+            �S@                          �5@�s.zqf@           P{@������������������������       ��T*E��?�            �s@������������������������       ���m�d@M            @_@                           @�)c���@�           �@                          �7@�i�"�@�           ��@������������������������       ��r�@�           ��@������������������������       �@��ɿ�@�            �r@                          �5@� i�[r@             ;@������������������������       �B8iY�o @             (@������������������������       ��:eϩ@             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     �s@     ��@     �@@     �J@     �}@     @R@     Џ@     �l@     �@     @v@      1@      $@     �k@     �s@      6@     �C@     �t@      M@     v@     �g@     �x@     `m@      .@      $@     `g@     �l@      5@      >@     �o@     �C@     `j@      a@     pq@      g@      *@      @     �b@     `h@      ,@      4@     �k@      ;@      h@     �\@      n@     �_@      *@             �F@     �Q@      @      @      E@      �?     �T@      8@     �[@     �A@       @      @     @Z@      _@      &@      0@     @f@      :@     �[@     �V@     @`@      W@      &@      @     �B@      B@      @      $@     �@@      (@      2@      7@     �C@     �L@              @      8@      0@      �?      �?      2@       @      @      .@      5@      >@              �?      *@      4@      @      "@      .@      @      &@       @      2@      ;@                      A@     �U@      �?      "@     @S@      3@     �a@      K@     �\@     �I@       @              2@      D@      �?      @     �@@      @     �M@      9@     �F@      .@      �?               @      :@      �?      @      $@      @     �E@      1@      ;@      @                      $@      ,@                      7@      �?      0@       @      2@      &@      �?              0@      G@              @      F@      ,@     �T@      =@     �Q@      B@      �?              �?      (@              �?      @      "@     �A@      @      4@      ,@      �?              .@      A@              @      D@      @      H@      7@      I@      6@                     �W@     �j@      &@      ,@     `b@      .@     Ȅ@      D@     0y@     @^@       @              .@     �T@      �?      �?     �A@      @     �q@      $@     �^@      8@       @                      1@      �?               @      @     �S@              9@      &@                              "@                      �?       @     �A@              &@      @                               @      �?              @      �?     �E@              ,@      @                      .@     �P@              �?      ;@      �?     �i@      $@     �X@      *@       @               @      J@              �?      .@              e@      @      K@      @       @              @      ,@                      (@      �?     �A@      @      F@       @                      T@     �`@      $@      *@      \@      &@     �w@      >@     �q@     @X@                      S@     ``@       @      &@     �Z@      $@     �w@      <@     0q@      X@                      K@     �[@      @      @     �N@       @     �s@      (@      g@     �P@                      6@      4@      @      @     �F@       @      P@      0@     �V@      =@                      @      �?       @       @      @      �?      @       @      @      �?                                               @      �?              @              @      �?                      @      �?       @              @      �?               @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJhl-,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@"�p@�	           ��@       	                    �?*�Z��@�           Ȗ@                          �0@+I}y@H           ��@                           �?�2R�~ @8            �T@������������������������       ���^�� @             7@������������������������       �X��v\A�?(             N@                           �?ȸ���H@           �{@������������������������       ��3Ǽ��@\            �c@������������������������       ����/*��?�            �q@
                            @�c��AN@9           �@                           �?�SЗ#}@�           ��@������������������������       ������@t             g@������������������������       �ظ�&�O@-           @~@                           �?�f��ݺ@�            `p@������������������������       ��� A�@             7@������������������������       ���ͥ?�@�            �m@                            @��'_�@!           .�@                            �?���Z@J           �@                          �8@w	���T@A           ��@������������������������       �HD?@           �@������������������������       �PhZ�2W	@&           �|@                           �?�t��	@	           �x@������������������������       �x�ٖ@E             Z@������������������������       ��c�j<�@�            @r@                          �=@�s�2	@�           ��@                           �?�-��Z	@�           �@������������������������       �E؀]O@g            �d@������������������������       ���}"@�	@:           �}@                          �?@�)����@6            @V@������������������������       ��>л�"@             J@������������������������       ����϶@            �B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@      p@     ��@      :@     �P@     `|@     �W@     �@     @m@     @�@      y@      ?@       @      O@      i@      @      $@     @a@      (@     @@     �S@     �s@     ``@       @              3@      L@                      D@       @     �m@       @     �`@      @@                      �?      3@                      (@              ?@              3@      �?                      �?      �?                      "@              @              @      �?                              2@                      @              8@              .@                              2@     �B@                      <@       @     �i@       @     �\@      ?@                       @      1@                      3@       @     �D@      @      E@      7@                      $@      4@                      "@             �d@       @      R@       @               @     �E@      b@      @      $@     �X@      $@     `p@     �Q@     �f@     �X@       @      �?      9@     @Y@      @      @      M@      @     �i@     �K@     `a@     @R@      �?      �?      ,@      :@               @      :@      @      :@     �@@      7@      ;@      �?              &@     �R@      @      �?      @@             @f@      6@      ]@      G@              �?      2@      F@       @      @      D@      @      M@      0@      F@      :@      �?      �?              @              @       @                      @      @       @                      2@      D@       @      @      C@      @      M@      $@      D@      8@      �?      *@     �h@     �v@      5@      L@     �s@     �T@     �~@     `c@     �|@     �p@      =@      &@     `a@     `o@      $@     �@@     `j@      K@     x@     �Y@     �t@     �f@      1@      "@     �[@     @h@      @      <@      c@      H@     �r@     �U@     �m@     �a@      ,@      �?      R@     �\@      @      2@      Y@      ;@      m@      B@      f@     �R@      @       @     �C@     �S@      �?      $@      J@      5@      P@      I@      O@      Q@      @       @      <@     �L@      @      @     �M@      @      V@      0@     �V@      C@      @               @      0@                      &@             �B@      �?      ;@      @               @      4@     �D@      @      @      H@      @     �I@      .@      P@      A@      @       @     �L@     �[@      &@      7@     @Z@      <@     @[@     �J@     @`@     �V@      (@      �?      K@     @W@      $@      1@     @U@      9@     �X@     �G@      _@      S@      (@              3@      =@              �?      2@             �C@      $@      D@      $@              �?     �A@      P@      $@      0@     �P@      9@      N@     �B@      U@     �P@      (@      �?      @      2@      �?      @      4@      @      $@      @      @      .@                              0@               @      $@      @      @      @              &@              �?      @       @      �?      @      $@              @       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�P_ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��z��W@�	           ��@       	                    �?>J��?Y	@           Ę@                          �<@{�q���@0           �~@                           �?!Kp��@           �z@������������������������       �yQZ0?Q@m            `e@������������������������       �����g�@�            p@                           �?�&w�@%            �N@������������������������       �����q@             B@������������������������       ��ex���@             9@
                           �?Q%V�	@�            �@                           �?��w@��@            z@������������������������       �ʐ�R�@d            �a@������������������������       ��V��	@�            @q@                           @*�Qz5
@�           @�@������������������������       �j��{h�	@�           P�@������������������������       ���{�Q	@;            �W@                           @߼����@�           0�@                          �=@��m+$�@�            �@                            �?�L@|�@l           ��@������������������������       �"sL���@�            Pt@������������������������       ���.��@�             o@                           @��\j�@             A@������������������������       �|�K-�@             5@������������������������       �W@���@             *@                          �4@{���@%           ��@                          �1@�P��A�@6           ��@������������������������       ���U���?�            �u@������������������������       �����1@`           ��@                          �6@ݷf��@�           0�@������������������������       ��;���@�            �r@������������������������       ��Jx��@7           �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �s@      �@      =@     �O@      |@     �T@     0�@     �i@     ؈@     `t@      A@      6@      g@     �n@      3@      @@     @n@     �J@     �k@     ``@     �n@      e@      5@             @P@     �V@      @      @     �P@      @     �Z@      ;@     �U@     �A@      �?              O@      S@      @             �I@      @     �Y@      6@      U@      6@      �?              *@      <@                      0@             @P@      @      B@      @      �?             �H@      H@      @             �A@      @      C@      1@      H@      .@                      @      ,@              @      .@              @      @      @      *@                      �?      *@              @      @               @      @      �?      @                       @      �?              �?       @              �?       @       @       @              6@     �]@     `c@      .@      ;@      f@      I@      ]@      Z@     �c@     �`@      4@      @      6@      P@      @      *@      R@      (@     �P@      B@      N@      M@      @       @      "@      @@               @     �C@       @      5@      @      .@      &@       @      @      *@      @@      @      &@     �@@      $@      G@      ?@     �F@     �G@       @      1@     @X@     �V@      (@      ,@      Z@      C@     �H@      Q@     �X@      S@      0@      ,@     @W@     @R@      $@      ,@     �V@      <@     �A@      L@     �W@     �P@      (@      @      @      2@       @              ,@      $@      ,@      (@      @      $@      @      �?     �`@     �r@      $@      ?@      j@      >@     p�@      S@     0�@     �c@      *@             �F@     �T@      �?      "@      S@      &@      f@      E@     �Z@      K@      @             �D@     @S@      �?      @      R@      @     �e@     �@@     �Z@      K@       @              8@     �C@      �?      @      E@      @      Y@      $@     @R@      7@       @              1@      C@                      >@      @     �R@      7@     �@@      ?@                      @      @               @      @      @      @      "@                       @              �?      @               @      @               @      @                       @              @      @                              @      �?       @                              �?     �V@     �k@      "@      6@     �`@      3@     �@      A@     �{@     �Y@      "@              B@     �Y@      @      (@      D@      @     �y@      0@      n@      H@       @              @      B@               @      &@             �f@      �?     �W@      .@       @              =@     �P@      @      $@      =@      @     �l@      .@      b@     �@@              �?      K@     @]@      @      $@      W@      0@     @l@      2@     �i@     �K@      @              @      N@      �?       @      C@       @     @V@             �T@      (@      @      �?     �I@     �L@      @       @      K@       @      a@      2@     �^@     �E@       @�t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?O���@�	           ��@       	                    @V��H�!@F           ��@                          �2@�*.���@           p�@                           �?	���3I@�            �p@������������������������       �3��&�@6            �T@������������������������       ����w9@o             g@                          �<@l���vI	@^           ��@������������������������       ��~�\�
	@           Љ@������������������������       ���LB�@W            �b@
                           @����S@C           ��@                            �?0
w���@           ��@������������������������       �?��@�            �t@������������������������       �����(@?           p~@                          �3@�٢�$@,             Q@������������������������       �y�'j��?             <@������������������������       �4a9��@             D@                          �5@C���@�           ԛ@                           @���\HZ@r           X�@                          �3@�<f�"C@K           @@������������������������       ��p�x|@�            �s@������������������������       �6��<:?@w            �g@                           @%8���@'           p}@������������������������       ���G��� @�            0v@������������������������       �݀اH@J             ]@                           @�@��@           P�@                           �?�W�4�a@N           �@������������������������       �ݣ�:�@N             \@������������������������       �;��G@            0y@                           �?������@�            pr@������������������������       �R�qԭ@8             U@������������������������       ����G�@�            `j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pq@     ��@      =@     �E@      z@      R@     Đ@      m@     h�@     pu@      =@      *@     �a@     �t@      *@      9@     �i@      H@     ��@     `a@      {@      i@      *@      *@     �\@     �g@      $@      2@     @b@     �E@     �k@     �[@     �k@      b@      (@       @      *@      G@                      ?@       @      U@      3@     �I@      2@      �?               @      @                      .@       @      5@       @      1@      $@      �?       @      &@      D@                      0@             �O@      &@      A@       @              &@     �Y@     �a@      $@      2@     �\@     �D@     @a@      W@     @e@     �_@      &@      "@      U@     �_@      $@      ,@     �Z@      ;@     �`@     @Q@      b@     �W@      "@       @      2@      1@              @      "@      ,@      @      7@      9@      @@       @              ;@      b@      @      @     �N@      @     `u@      <@     �j@     �L@      �?              7@     @`@       @      @      N@      @     pt@      7@     `i@      D@      �?              $@      F@      �?              9@      �?     �b@      $@      R@      4@                      *@     �U@      �?      @     �A@      @      f@      *@     ``@      4@      �?              @      ,@      �?      �?      �?              .@      @      $@      1@                              @              �?      �?              &@              �?      $@                      @      $@      �?                              @      @      "@      @              @     �`@     �p@      0@      2@     `j@      8@     �@     @W@     �u@     �a@      0@      @     �G@      a@      @      @     @X@      1@     v@      I@     �g@     �L@       @      @      ?@      S@      @       @     �R@      $@      _@     �C@      W@      D@      @       @      9@     �A@              �?     �F@      @     �V@      8@     �I@      A@       @       @      @     �D@      @      �?      =@      @      A@      .@     �D@      @      @              0@      N@      �?      @      7@      @     �l@      &@     �X@      1@      @              *@     �F@              @      .@       @     �g@      @      Q@      &@                      @      .@      �?      �?       @      @     �C@      @      ?@      @      @      �?      V@      `@      (@      &@     �\@      @     �c@     �E@     �c@     @U@       @      �?     @R@      W@       @      @     �R@      @     �Q@     �A@      S@      P@       @              ,@      (@      @      @      3@              <@      @      &@      2@      �?      �?     �M@      T@      @      @      L@      @      E@      @@     @P@      G@      @              .@     �B@      @      @     �C@      �?     �U@       @      T@      5@                      @      *@                      @              >@              9@      @                      (@      8@      @      @      @@      �?      L@       @     �K@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���XhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @M�+ؼ�@�	           ��@       	                   �3@��/��@m           B�@                           @����R�@�           @�@                          �1@hQ^Ƥ�@c            �@������������������������       �^FW�>@�             k@������������������������       �X!h@�            �v@                           @&4�Y@Y            �`@������������������������       �ש*���@P             ^@������������������������       �]<����@	             (@
                          �<@_M���q	@�           d�@                           �?���֭>	@           T�@������������������������       �ud�~�t	@K           @�@������������������������       �J/L_ɛ@�            �r@                           �?D�
��@�            @p@������������������������       �,���,@$             M@������������������������       �`�Q�@v            @i@                           �?���,�h@           ��@                           @�<����@[           ��@                          �4@��q`3� @�            `v@������������������������       �;�v����?�            �n@������������������������       �t��䃾@C            �\@                            �?;�l���@�            �i@������������������������       �<!�;|��?            �C@������������������������       ���:m �@d            �d@                           @��xΐd@�           ؑ@                           @��~��@�           ��@������������������������       �=L\
@�            �p@������������������������       �����Í@W           0�@                           �?iEe�:@�            `t@������������������������       ����$�( @             8@������������������������       ��iͱ�9@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     Ps@     x�@      9@      L@     �{@      W@     x�@      o@     ��@      x@      :@      4@      l@     �s@      .@      C@     @s@     @Q@     �v@     �j@     v@     �p@      6@      @      F@      W@       @      @     @V@      .@      g@      K@      b@     �S@      �?             �B@     �Q@       @      @     @R@      @      d@      @@     �_@     �P@                      "@      ;@       @      �?      2@             �S@      ,@     �J@      .@                      <@      F@              @     �K@      @     �T@      2@     �R@     �I@              @      @      5@                      0@       @      7@      6@      2@      (@      �?      @      @      4@                      (@      @      7@      6@      0@      (@              �?              �?                      @      @                       @              �?      0@     �f@     �k@      *@      A@     `k@      K@     �f@      d@      j@     �g@      5@      (@     �b@     `f@      &@      ;@     @g@     �@@      e@     �_@     �g@     �`@      4@      (@     ``@     �`@      $@      4@      a@      8@      Y@      Y@     @b@     �Z@      3@              3@     �G@      �?      @      I@      "@      Q@      :@     �F@      <@      �?      @      ?@     �D@       @      @     �@@      5@      ,@      A@      1@     �K@      �?              "@      $@      �?      �?      @      @      @      @       @      0@              @      6@      ?@      �?      @      =@      0@      @      ?@      .@     �C@      �?       @      U@     �n@      $@      2@     `a@      7@     �@     �A@     �y@     �]@      @              2@     �T@       @       @      =@      @      p@      "@     @`@      ;@      �?              *@      L@                      ,@      @      f@      @      S@      (@                      &@      :@                      @             �`@      �?      K@      $@                       @      >@                      @      @     �D@      @      6@       @                      @      ;@       @       @      .@              T@      @      K@      .@      �?                      �?       @              @              3@              $@                              @      :@               @       @             �N@      @      F@      .@      �?       @     �P@     �d@       @      0@     �[@      2@     v@      :@     �q@      W@      @       @      F@     �_@      �?      @     �N@       @     r@      1@     �h@     @P@      @       @      3@      L@              �?      <@       @     @S@       @      H@      0@      @              9@     �Q@      �?       @     �@@             �j@      "@     �b@     �H@                      6@      C@      @      *@     �H@      $@      P@      "@     �U@      ;@                      �?                              @              �?      @      &@      �?                      5@      C@      @      *@     �E@      $@     �O@      @      S@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJd�[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�6PB>@�	           ��@       	                    �?(���@�           �@                           �?E0���^@3           ��@                            �?Q8�b@            |@������������������������       ��ǀ)�@�            �t@������������������������       �L-��@J            �]@                          �5@�Lo ��@           0{@������������������������       ��ǿ?MJ@�            �p@������������������������       �$���oM@l             e@
                          �4@���=�@�           �@                          �3@S��>@%           �@������������������������       ���d\�@�           H�@������������������������       �Ϯ���@�             k@                           @A�D��@�           �@������������������������       ��v�v�	@a           �@������������������������       ��q�kU@*           P~@                           @!�Y�@�           L�@                           �?1�O:��@&           ��@                          �6@uz����@�            �o@������������������������       ��a�@~@^            �b@������������������������       �@��x��@>            �Y@                           �?K@eV�q	@�           ��@������������������������       ����$�	@�             j@������������������������       ���G��@�            `x@                           �?b��np�@�            p@                           �?3/`1���?5            �T@������������������������       ��B/���?            �E@������������������������       � �M]�x�?             D@                          �1@OԲY@r            �e@������������������������       ��t���)�?             :@������������������������       ���	@c            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     t@     ȁ@      ?@      K@     �{@      V@     ��@     �h@     p�@     �u@      :@      &@     �k@     �x@      (@      D@     s@      K@     ��@     �a@     Ѓ@     �n@      1@      �?      L@      a@      @      @     �Q@      $@     �s@      :@      i@      K@      @      �?      ;@     �Q@      �?      @     �B@      @     �f@      *@      S@      >@      �?      �?      5@      H@      �?      @      @@      @      `@      (@     �I@      :@      �?              @      7@                      @       @      J@      �?      9@      @                      =@     @P@       @             �@@      @     `a@      *@     @_@      8@       @              .@     �D@                      @             �Z@      @     �S@      .@                      ,@      8@       @              ;@      @     �@@       @      G@      "@       @      $@     �d@      p@      "@      B@     `m@      F@     �y@     �\@     {@      h@      ,@             �N@     @_@      @      (@     �W@      (@     pp@     �A@      i@      U@      @              E@     �W@      @      &@      M@      &@     �j@      <@     `d@      L@      @              3@      ?@      �?      �?      B@      �?     �I@      @     �B@      <@      @      $@      Z@     ``@      @      8@     �a@      @@      c@     �S@      m@      [@      @      "@     @P@      S@      @      2@     �R@      8@     �G@     �N@      X@      O@      @      �?     �C@     �K@       @      @     �P@       @     @Z@      2@      a@      G@       @      @      Y@      f@      3@      ,@     `a@      A@     @n@     �L@     �j@     �X@      "@      @     �V@     �a@      .@      ,@     @]@     �@@     �b@     �L@      a@     �T@      @              <@      G@      @      @      @@      @      O@      "@      H@      .@                      1@      >@              �?      (@      @     �H@       @      ;@       @                      &@      0@      @      @      4@              *@      @      5@      @              @     �O@     @X@      (@       @     @U@      >@     �U@      H@      V@      Q@      @       @      5@      B@      $@      @      ?@      (@      :@      "@      ;@      <@       @      @      E@     �N@       @      @      K@      2@      N@     �C@     �N@      D@      @              "@      A@      @              6@      �?     �W@              S@      .@       @              �?      @                      @              E@              ?@      �?                      �?      @                      �?              7@              ,@      �?                               @                       @              3@              1@                               @      =@      @              3@      �?      J@             �F@      ,@       @                      @                                      3@               @                               @      8@      @              3@      �?     �@@             �E@      ,@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�(QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?&J�JM@�	           ��@       	                    �?��X�Uk@           ԓ@                           �?$����@*           �~@                            �?\,�g@�@o            @f@������������������������       ��|
��@            �H@������������������������       ��,7�@S             `@                            @��՚Uh@�            �s@������������������������       �|��/�8@c            �c@������������������������       �z+;���@X            �c@
                          �4@֠�_m2@�           H�@                           @����� @!           0|@������������������������       �ØS�{@:            @W@������������������������       ��o꘹w�?�            `v@                          �7@
�7e�@�            `t@������������������������       �bX<��@j            �d@������������������������       ���c:O@h            �c@                           @�SX�M@�           ��@                          �7@놁a'@U           �@                          �3@5��,�-@H           <�@������������������������       �ە�`"�@            �@������������������������       �Jqw.@/           X�@                           �?eƴ��I	@           Љ@������������������������       ��Wǈ0I	@4            �T@������������������������       ���u�	@�           8�@                          �4@��Q�@	@0            �R@                            @���JF�@             9@������������������������       ��GE��� @	             .@������������������������       ����N�@             $@                           �?��0�*�@              I@������������������������       �/p3O�@	             .@������������������������       �h��%1@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      q@     �@      ?@     �P@     �|@     @T@     l�@     �i@     �@     x@      @@             @S@     �c@      @      "@     �\@      $@     0}@      H@     �q@     �V@      @             �I@     @R@      �?      @     @Q@      @     @\@      <@     @X@      I@                      0@      0@                      8@             �L@      @      H@      *@                       @      @                       @              (@       @      3@      @                      ,@      *@                      0@             �F@       @      =@      $@                     �A@     �L@      �?      @     �F@      @      L@      8@     �H@     �B@                      2@      :@      �?      �?      ,@      @      ;@      &@     �@@      5@                      1@      ?@              @      ?@       @      =@      *@      0@      0@                      :@     �U@      @      @      G@      @      v@      4@     �g@      D@      @              5@      C@              @      ,@             �m@      &@     @Z@      4@      �?               @      @               @      @              =@      @      @@      @                      *@     �@@              @       @             �i@      @     @R@      *@      �?              @      H@      @              @@      @     �]@      "@     @U@      4@       @               @      @@      @              9@       @     @Q@      �?      >@      @                      @      0@                      @       @     �H@       @     �K@      1@       @      2@     �h@      x@      ;@     �L@     �u@     �Q@     @�@     �c@     �}@     pr@      =@      *@      g@     �w@      ;@      L@     �t@      P@      �@     �b@     @}@      r@      <@      @      a@     �p@      "@      D@     �h@      :@     �}@     @T@     0t@     `d@      0@      @     �D@      _@       @      $@     �S@      &@     �q@      E@      e@     �W@      @      @     �W@     `b@      @      >@      ^@      .@      g@     �C@     @c@      Q@      (@      @     �H@     �[@      2@      0@      `@      C@      [@     �Q@      b@     @_@      (@      @      @      @              @      1@      @       @       @      (@      0@      @      @      E@      Z@      2@      &@      \@      A@     �Z@      O@     �`@     @[@      "@      @      (@      @              �?      0@      @      @      @      $@      @      �?              @       @              �?      �?      �?      @      �?      @      @      �?              @                      �?                      �?      �?      �?      @                               @                      �?      �?       @              @              �?      @      @      @                      .@      @      �?      @      @      �?              @                                      @      @      �?      �?              �?               @      @      @                      "@      @              @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�9�q7A@�	           ��@       	                    �?΍�V?@�           ��@                          �8@t4��@�            0t@                           �?���@�             p@������������������������       ��7����@;            �U@������������������������       ��(���M�?i            �e@                           �?7�Yq�S@(            @P@������������������������       ��41X�@             A@������������������������       ������@             ?@
                           @MGds�@�           ȅ@                           �?�L<��9	@           �{@������������������������       ��"���@Q            �`@������������������������       �&����~	@�            �s@                          �1@�Bil�@�            `o@������������������������       �W	p��?            �C@������������������������       ��[��<@�            �j@                           @�ރ�E@5           ��@                          �1@;���f�@�           t�@                           @6��X@o            �f@������������������������       �������@T            @a@������������������������       �N�ɫ@             F@                           �?�
�& 	@_           ��@������������������������       ��1-��n	@�           ��@������������������������       ��DI�Tm@�             u@                           �? u���@g           ��@                           @>g��Q@           �|@������������������������       ����S��?�            �m@������������������������       ��H�{@�             l@                          �7@A�� @J           �@������������������������       �Ѵ� ��@�           ��@������������������������       ��+x\C@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      r@     P�@      @@     �I@     �|@     @W@     @�@      j@     ��@     �u@      =@      @     �T@     @`@      @      *@      ]@     �@@     pr@      M@     �i@     �P@      *@      @      ,@      B@               @      @@      @      `@      @      T@      ,@      @               @      9@               @      @@      �?     @\@      @      P@       @      �?              @      (@              �?      &@              5@      @      :@      @      �?              �?      *@              �?      5@      �?      W@              C@      @              @      @      &@                              @      .@      �?      0@      @       @      @      @      @                              �?       @      �?      @      @                       @      @                              @      @              "@      @       @              Q@     �W@      @      &@      U@      ;@     �d@     �J@     �_@     �J@      $@             �F@      P@       @      $@      P@      9@     �P@     �H@     �O@     �G@      $@               @      3@              @      ,@       @      >@      ,@      ?@      "@      �?             �B@     �F@       @      @      I@      7@     �B@     �A@      @@      C@      "@              7@      >@       @      �?      4@       @      Y@      @     �O@      @                              @              �?      �?              <@      �?      @       @                      7@      ;@       @              3@       @      R@      @      N@      @              1@     �i@     �z@      <@      C@     �u@      N@     H�@     �b@     H�@     pq@      0@      .@     @b@     @m@      3@      ;@     �k@     �E@     @m@      _@      l@     �i@      $@      @      @     �B@      �?              4@              J@      *@      @@      3@                      @      ;@      �?              1@             �G@      @      :@      "@              @      �?      $@                      @              @      @      @      $@              (@     �a@     �h@      2@      ;@      i@     �E@     �f@     �[@      h@      g@      $@      (@     �Z@     �b@      .@      9@      c@     �A@      [@     �S@     `a@     �b@      $@              A@     �H@      @       @     �G@       @     �R@      @@      K@     �A@               @      N@     �g@      "@      &@      _@      1@     �@      ;@     �v@     �R@      @              2@     �O@               @      9@      @      k@      @     �[@      2@                      *@      =@                      "@      @      `@       @     �G@      @                      @      A@               @      0@              V@      @     �O@      *@               @      E@     �_@      "@      "@     �X@      *@     pr@      5@     @o@     �L@      @              6@     �Y@      @      @     �J@      *@     �n@      $@     �h@      B@      @       @      4@      9@       @       @      G@              I@      &@     �I@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ�lvhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?)�Ǒ@�	           ��@       	                   �8@:$H�@�           X�@                           �?94��@�           �@                          �5@p��e�@�             r@������������������������       ���;� @}            @i@������������������������       ���&�WU@2             V@                           @A�a�@J           ؀@������������������������       ��#���@�            �l@������������������������       �n�}���@�            ps@
                          �<@H�eN	@�            �q@                           �?4#����@r            �e@������������������������       ��{,jѐ@6            �U@������������������������       ��+��n@<             V@                           @A��V<�@?            �Z@������������������������       �ͽ��t	@/            �S@������������������������       �E�����@             =@                           �?qk�fF�@�           �@                           �?�龝?�@�           ̑@                            @R�Y��@�            `v@������������������������       ��ㅩL�@d            �c@������������������������       �g� h>@|             i@                          �:@��r�f	@�           h�@������������������������       �S%!	@�            �@������������������������       ���m	@^            �a@                           @�t�w�@.            �@                           �?�z>|�@�           ��@������������������������       �G����v@�            `l@������������������������       �2D�@-           �}@                          �1@�;�3�@v           �@������������������������       �v�����?             i@������������������������       �z��f@�           ȇ@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@     ȁ@      7@      L@     0~@     �S@     T�@     �g@     ��@     `u@      =@      @     �W@     �b@      @      2@     �b@      8@     Ps@      O@      i@      U@      (@             @S@     �]@       @      (@      ]@      &@     �p@      A@      c@     �E@                      (@      E@      �?      @      :@      �?      `@       @     @P@      "@                      @      <@              @       @      �?     �V@       @      M@      @                       @      ,@      �?      �?      2@             �B@              @       @                     @P@      S@      �?       @     �V@      $@      a@      @@     �U@      A@                     �A@      3@               @     �H@       @      N@      &@      >@      4@                      >@     �L@      �?      @     �D@       @      S@      5@     �L@      ,@              @      2@     �@@      �?      @      @@      *@     �F@      <@     �H@     �D@      (@      @      *@      8@      �?       @      1@      @     �B@      3@     �A@      .@      @      �?      @      ,@      �?       @      @      �?      1@      $@      2@       @      @       @      "@      $@                      &@      @      4@      "@      1@      @                      @      "@              @      .@      "@       @      "@      ,@      :@       @              @      "@              @      *@      @       @      @      &@      *@      @                                               @       @              @      @      *@      @      *@     `i@      z@      4@      C@     �t@     �K@      �@     �_@     8�@      p@      1@      (@     �Z@     `i@      .@      0@     �e@     �A@      g@     �Q@      c@     �c@      .@              >@     @P@      �?      @      K@      @     �S@      1@     �O@      C@       @              .@      5@      �?       @      :@              <@      @      A@      8@       @              .@      F@              @      <@      @     �I@      (@      =@      ,@              (@      S@     @a@      ,@      &@     �]@      ?@     @Z@      K@     @V@     �]@      *@      @      M@     �^@      $@      @      W@      9@     �X@      F@      S@     @V@      (@      @      2@      0@      @      @      ;@      @      @      $@      *@      >@      �?      �?     @X@     �j@      @      6@     @d@      4@     @�@      L@     �z@     @Y@       @      �?     �K@     �X@      �?       @     @T@      2@      i@      >@     �d@      E@      �?              0@      =@                      3@       @     �W@      @     �K@      @              �?     �C@     �Q@      �?       @      O@      0@     �Z@      8@     �[@      B@      �?              E@      ]@      @      ,@     @T@       @     �u@      :@     �p@     �M@      �?              "@      ,@                      ,@              [@             �H@      @                     �@@     �Y@      @      ,@     �P@       @     `n@      :@      k@     �J@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-��vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Y+�X�z@�	           ��@       	                    �?�!�	@[           ��@                           �?¶=��	@�           ��@                           �?3�@w�`@�           �@������������������������       �����Ӷ@�            �p@������������������������       ��g"���@�            pw@                           �?z�j��	@i           ��@������������������������       �t�ђ�@�            �p@������������������������       ��[}Fsn
@�           ��@
                           �?��2�@@r           Ђ@                            �?~�
vŽ@m            `e@������������������������       ���gՈF @%             M@������������������������       ��]��+@H            @\@                          �3@�	-�@           �z@������������������������       ����@@c            �d@������������������������       ��C\�c�@�            �p@                          �7@QSU 0@@           8�@                           �?�̔��@7           ��@                           @�������?)           `~@������������������������       �M܏ȡ@�?�            `u@������������������������       �L��Ζ�@W             b@                           @��1b{M@           @�@������������������������       �g�k8��@p            �g@������������������������       �e[ٷu�@�           P�@                            @��"R@	            z@                           @��|o0�@�            �t@������������������������       �;�z3@�            �j@������������������������       �������@N            �^@                           �?8<A#��@2            @T@������������������������       ������?            �@@������������������������       ���F%��@             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     `q@     8�@     �A@     �Q@     �z@     �S@     ��@      m@     �@     Pv@     �C@      4@     `i@     �s@      8@      K@     `r@      N@     �v@     �f@     Pw@     �n@      =@      4@     �b@     �k@      4@     �E@      k@      F@     �m@     �b@     �n@      h@      <@      @     �A@     @W@      @      ,@      V@      "@     �`@      M@     �[@     �R@      ,@      @      1@     �F@      @      @      F@      @      I@      1@     �F@      9@      @      �?      2@      H@      �?      "@      F@      @     @U@     �D@     �P@      I@      @      ,@      ]@      `@      0@      =@      `@     �A@     �Y@     @W@     �`@     @]@      ,@              >@     �D@      �?      @      @@      @      H@      9@      H@      @@      �?      ,@     �U@     �U@      .@      6@     @X@      @@      K@      Q@     �U@     @U@      *@              J@     @X@      @      &@     @S@      0@     @`@      @@      `@      K@      �?              1@      2@                      6@      �?      K@      @     �G@       @                       @      $@                       @      �?      4@              6@      �?                      .@       @                      4@              A@      @      9@      @                     �A@     �S@      @      &@     �K@      .@      S@      <@     @T@      G@      �?              &@      7@              �?      2@       @     �I@      @     �A@      1@                      8@      L@      @      $@     �B@      *@      9@      5@      G@      =@      �?      �?     �R@      m@      &@      1@     �`@      2@     h�@     �H@     �z@     �[@      $@             �J@      i@       @      *@     �S@      &@     (�@      ,@     �s@     �Q@      "@              &@     @P@              @      3@      �?     0p@       @     �Y@      2@      �?              $@     �E@                      &@      �?      h@      �?     �R@      $@                      �?      6@              @       @             �P@      �?      =@       @      �?              E@      a@       @      @      N@      $@      r@      (@      k@      J@       @              ,@     �D@                      (@      @      O@      @      >@      *@      @              <@     �W@       @      @      H@      @     �l@      @     @g@     �C@       @      �?      6@      @@      @      @     �K@      @      Z@     �A@     �[@     �D@      �?      �?      4@      >@       @       @      H@      @     �Q@      =@     �V@     �A@      �?      �?      &@      7@                      A@      �?     �J@      (@      M@      2@      �?              "@      @       @       @      ,@      @      1@      1@      @@      1@                       @       @      �?       @      @              A@      @      5@      @                              �?              �?                      3@       @      "@      �?                       @      �?      �?      �?      @              .@      @      (@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJÕ�WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?V�h�Au@�	           ��@       	                     @�0s���@           l�@                          �4@��
��@?           h�@                           @W�i@3           p~@������������������������       �\��\;j@t            �f@������������������������       �{{�W� @�             s@                           �?��5_"'@           `z@������������������������       ��=�o@�            �k@������������������������       �PE�0�@�            @i@
                           @���_�+@�            �t@                          �8@kΐ��h@�            �n@������������������������       ����_�)@v            �e@������������������������       �0�R\��@-            �Q@                           @N�۾C��?6             V@������������������������       ��#OK |�?             D@������������������������       ��x^2�$�?              H@                          �5@Y�t+�L@�           ܤ@                           @���2k�@l           ԕ@                           �?rD�F�@�           ��@������������������������       ����ߟ6	@6            @������������������������       �7��͙�@�            �m@                           @�D�,D�@�           ��@������������������������       ���[5�6@�           @�@������������������������       �jg���@	             .@                           @T��`G&	@           �@                          �8@Q+��I�	@�           �@������������������������       �c��e@�            �u@������������������������       ��bǺ��	@           p|@                          �6@b����@#           �}@������������������������       ��HMH@=            �X@������������������������       ����{�@�            Pw@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     ��@      8@     �Q@     }@     @X@     ��@     �k@     �@     �t@      9@              Z@      f@      @      ,@     �\@      &@     pz@     �E@     �q@     @Q@      @             �Q@     `a@       @      @     �S@      &@     �s@      9@     `i@     �J@      @              8@     �O@              @      =@             �j@      $@     @\@      <@       @              .@      >@               @      ,@             �J@      @      H@      0@                      "@     �@@              @      .@              d@      @     @P@      (@       @              G@      S@       @              I@      &@      Z@      .@     �V@      9@      @              <@      A@      �?              8@       @     @P@      "@     �A@      0@                      2@      E@      �?              :@      @     �C@      @     �K@      "@      @              A@     �B@      �?      "@     �A@             �Z@      2@     �S@      0@                      @@      A@      �?      @      ?@              L@      0@      K@      .@                      0@      5@      �?       @      6@             �I@       @     �E@      &@                      0@      *@              @      "@              @       @      &@      @                       @      @               @      @              I@       @      8@      �?                      �?      @                                      ;@              "@                              �?                       @      @              7@       @      .@      �?              5@     �j@      x@      5@      L@     �u@     �U@     p�@     @f@     P�@     Pp@      4@      &@      P@     `i@       @      =@     @c@     �A@     @w@      R@     �t@     �[@      "@      &@      B@     �[@      @      0@     �\@      9@     `a@      P@     @`@     �S@      @      &@      @@     �O@      @      .@     @U@      3@      S@      C@     �V@     �M@      @              @     �G@       @      �?      =@      @     �O@      :@     �C@      3@                      <@     @W@      @      *@      D@      $@      m@       @      i@      @@      @              <@     �V@      @      (@     �C@      @      m@       @     �h@      =@      @                       @              �?      �?      @                      @      @              $@     �b@     �f@      *@      ;@     �h@     �I@     @g@     �Z@      h@     �b@      &@      "@     �X@      _@      @      7@     �_@     �E@     �Q@     �U@      V@     �\@      &@       @     �H@      P@      @      ,@      S@      "@      4@      4@      F@     �D@      @      @     �H@      N@      @      "@     �I@      A@     �I@     �P@      F@     @R@      @      �?      I@     �L@      @      @     �Q@       @     �\@      4@      Z@     �B@                      *@      "@      @              0@             �D@              (@      @              �?     �B@      H@      @      @      K@       @     �R@      4@      W@      @@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�)<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @)�-YA^@�	           ��@       	                    �?�����@p           ġ@                          �<@r�O�]@�           ��@                           �?��C�W@i           x�@������������������������       �xp�}r@	           P{@������������������������       �ل��c @`            @c@                            �?֝�`�@-            @Q@������������������������       ��r�-�@            �I@������������������������       � l\�o�@             2@
                          �1@�!/q;U	@�           8�@                           @��F��@d             d@������������������������       ��3�`�@[            @b@������������������������       �^,Eal�@	             ,@                          �9@�+���	@v           ��@������������������������       ��s��	@z           L�@������������������������       �9���	@�            �y@                          �6@+��a�=@           ��@                          �1@e�G��@�           �@                           @��8E�* @�            �s@������������������������       �\	�v��?�            �l@������������������������       ��P��=@5            �U@                           �?m}u��@           X�@������������������������       �7`��<@ @�            @p@������������������������       ���
�$@d           8�@                            @��!"�@2           ~@                           �?XN2���@�            �x@������������������������       �R�e(�@�            `j@������������������������       ���yA@w            @g@                           @2?5Ľ�@6             U@������������������������       ���%���?             D@������������������������       ��S1&�@             F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     ��@      @@      J@     �|@     �R@     h�@     �j@     ��@     @w@     �A@      2@     �j@     �u@      6@      C@     0s@     �N@     `x@     �f@      y@     �p@      >@       @      Q@      U@       @       @     @Q@      @     @f@      5@     �c@     �O@      @       @     �N@     �Q@       @      @      O@      @     �e@      1@     �b@      E@      @       @     �H@     �O@       @      @     �I@      @      [@      1@     @Y@      A@      @              (@       @                      &@             �P@              H@       @                      @      *@              @      @              @      @       @      5@       @              @      @              �?      @              �?      @      @      5@       @              �?      @              @       @               @      �?       @                      0@     @b@     `p@      4@      >@     �m@      M@     �j@     �c@     �n@     `i@      9@              &@      ;@      �?              &@       @     �F@      2@      D@      @                      $@      ;@      �?              @              F@      0@     �B@      @                      �?                              @       @      �?       @      @                      0@     �`@     `m@      3@      >@     `l@      L@     �d@     �a@     �i@     �h@      9@      $@      V@     `f@      ,@      6@     �g@      8@      a@      V@     @b@      `@      1@      @     �G@      L@      @       @      C@      @@      >@     �J@     �M@     @Q@       @      @     �T@     @k@      $@      ,@     �c@      *@     8�@     �@@     �y@     �Z@      @              K@     �c@      @      "@     @W@      @     p}@      *@     `q@     @P@      @              (@      7@              @      1@             �c@      �?     @U@      2@                       @      (@                      $@              `@             �L@      *@                      @      &@              @      @              <@      �?      <@      @                      E@     �`@      @      @      S@      @     �s@      (@      h@     �G@      @               @      G@               @      ,@              `@       @      K@      @                      A@      V@      @      @      O@      @     `g@      $@     `a@     �D@      @      @      =@     �N@      @      @     �O@      @      \@      4@      a@     �D@      �?      @      ;@      M@      �?       @     �L@      @      T@      0@      ]@      @@      �?      @      6@      B@               @      ;@      �?     �D@       @     �I@      3@      �?              @      6@      �?              >@      @     �C@       @     @P@      *@                       @      @       @      @      @       @      @@      @      5@      "@                       @                               @       @      4@              *@      �?                              @       @      @      @              (@      @       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@]�K�\@�	           ��@       	                   �2@f��Je�@           .�@                           @z��L��@�           ��@                           @�4�y�@$           �|@������������������������       �����7�@�            �w@������������������������       �}�7�_�@3            �S@                            �?��(�� @a           8�@������������������������       �0�w���?K             _@������������������������       �	���@           �z@
                           @.�d��@�           ��@                           �?� ��E@N           ��@������������������������       �;`��d�@`           �@������������������������       ��t+�@�            �w@                           @
	Y�I]@9           �~@������������������������       ���&�?l            �f@������������������������       ��T�@�            0s@                           �?}%X�	@�           Ȗ@                          �8@o4r�"�	@�           P�@                            �?@p�Ga@�            �k@������������������������       �	��%q@A            @[@������������������������       ����)�|@K            @\@                           �?����	@N           `�@������������������������       �hbeI�@p            �f@������������������������       �Vq�ʾ�	@�            pw@                           @���-r@�           @�@                            @ե*m�@�            @j@������������������������       ��4�1��@]             b@������������������������       �O	N��@(            �P@                          �<@��k��d@4           `}@������������������������       ��4cCg�@�            �w@������������������������       �́L^e@7            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     ��@      <@     �F@     `}@     �W@     ��@     �k@     ��@     �u@     �B@      &@     �b@     �v@      ,@      2@     `p@      A@     X�@      Z@     x�@     `f@      ,@      @     �D@     �`@      �?      @     �Y@      @     �y@      F@     �i@     �L@      �?      @      9@     �P@      �?      �?      O@      @      b@     �@@     �R@     �D@      �?       @      3@      E@      �?      �?      J@      �?     �`@      7@      R@     �A@               @      @      9@                      $@       @      *@      $@      @      @      �?              0@     �P@              @     �D@             �p@      &@      `@      0@                       @      1@                      @             �S@              2@      @                      ,@      I@              @      B@             �g@      &@     �[@      *@              @      [@     �l@      *@      *@     �c@      ?@     �v@      N@     0t@     �^@      *@      @      X@      e@      $@      $@     @[@      =@     �d@      L@     �h@      X@      (@      @     @P@     �Y@      @      @     �R@      1@     @Q@     �C@      \@     @Q@      (@              ?@     �P@      @      @      A@      (@     @X@      1@      U@      ;@                      (@     �N@      @      @      I@       @      i@      @     �_@      :@      �?              @       @                      1@             �V@      @     �L@      @                      "@     �J@      @      @     �@@       @     �[@      �?     �Q@      5@      �?      @     �b@      i@      ,@      ;@      j@      N@     `j@      ]@     �p@     `e@      7@      @     �V@     �Y@      &@      3@      `@     �C@     �T@     �Q@     @Y@      Z@      7@              :@      @@      @      $@     �H@      @      7@      "@      F@      .@      @              .@      "@      @      @      8@       @      "@      @      9@      @       @              &@      7@       @      @      9@      �?      ,@       @      3@      $@      @      @      P@     �Q@      @      "@      T@      B@     �M@      O@     �L@     @V@      2@      @      *@      :@              �?      @@      @      ?@      *@      4@      =@       @      @     �I@     �F@      @       @      H@      ?@      <@     �H@     �B@      N@      $@              N@     �X@      @       @     �S@      5@      `@     �F@     @e@     �P@                      <@      A@              @      9@      @      ?@      5@      B@      :@                      *@      3@              @      7@      @      1@      &@      @@      4@                      .@      .@                       @              ,@      $@      @      @                      @@      P@      @      @      K@      0@     �X@      8@     �`@     �D@                      5@      K@      �?      @      A@      (@      V@      7@     �\@      =@                      &@      $@       @      �?      4@      @      $@      �?      4@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�q hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��h@�	           ��@       	                    �?��͍��@           ��@                            �?�C�JM@-           0@                           �?����a�@N            @a@������������������������       �8ՒA҅@$            �P@������������������������       � ���@*             R@                            @�}��P@�            �v@������������������������       ����Ɨ@`            @b@������������������������       �'XJkd@            �j@
                          �>@u8M$>+@�           ��@                          �3@�t�&�� @�           �@������������������������       �0a����?�            �v@������������������������       ����P�@�            `w@������������������������       ����v�t@             ,@                           �?W����@�           ʤ@                            @����2O	@�           $�@                          �<@-?��~X	@�           ��@������������������������       ��/Ks�I	@s           0�@������������������������       ���Q[0�@2            �R@                           @�U<�	@&           �}@������������������������       �-Wc�j�@           `z@������������������������       �`�1Ó@             I@                           �?���[E@�           p�@                           @���Dg@9            �X@������������������������       �^,\�@            �F@������������������������       �DIS�]9@!             K@                           @��`�@�           �@������������������������       ���jm��@           �@������������������������       ��M�=^@x            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        &@     �r@     ��@      ;@      O@     �z@     �S@     ,�@     �j@     ��@     �w@      5@      �?     �R@     @f@      @      "@     @X@      @     �~@      D@     �p@     �S@       @      �?     �I@      U@       @      @     �N@              ^@      6@     �Y@      G@       @      �?      (@      ?@                      3@              <@      @      >@      $@      �?      �?       @      *@                      $@              5@      @      &@      @                      $@      2@                      "@              @       @      3@      @      �?             �C@     �J@       @      @      E@              W@      0@     @R@      B@      �?              $@      ,@      �?       @      3@              D@      @      C@      .@      �?              =@     �C@      �?      @      7@              J@      $@     �A@      5@                      8@     �W@       @       @      B@      @     pw@      2@     �d@      @@                      8@     �W@       @       @     �@@      @     pw@      ,@     `d@      <@                      .@      >@                      "@              i@       @     �V@      &@                      "@      P@       @       @      8@      @     �e@      @      R@      1@                                                      @       @              @      �?      @              $@     @l@     �v@      7@     �J@     �t@     @R@     ��@     �e@     8�@     �r@      3@      "@     �^@     `c@      *@      6@     �f@      E@     �Z@      [@      e@     `c@      0@      @     �P@     �U@      @      ,@      W@      8@     �P@     @S@      U@     �W@       @      @     �L@     �T@      @      *@     �S@      3@     �P@     �P@     �S@     @R@      @      �?      $@      @              �?      *@      @              &@      @      6@       @      @     �K@      Q@      @       @     @V@      2@      D@      ?@      U@      N@       @      @      K@     �L@      @       @     �S@      1@     �A@      =@     @S@     �I@      @      �?      �?      &@                      $@      �?      @       @      @      "@      @      �?      Z@      j@      $@      ?@     �b@      ?@      {@     @P@     �w@     �a@      @      �?      @      ,@              (@      @      @      *@      "@      7@      &@              �?      �?       @              &@      @      @      �?      @      �?       @                      @      @              �?      �?              (@      @      6@      @                     �X@     `h@      $@      3@     �a@      ;@     Pz@      L@     �v@     �`@      @             �R@     �e@      $@      1@     @_@      4@     0w@      F@     �t@     @[@      �?              9@      6@               @      2@      @      I@      (@      >@      7@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJyV
.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�jh~8@�	           ��@       	                    �?�ьGs�@i           �@                            �?zI�-�:@�           @�@                           �?Ll�6/@u            @g@������������������������       ���P~�@9            �V@������������������������       �D�� �@<             X@                           �?N;�b@           �z@������������������������       �k�I�!@�            �r@������������������������       ��]#2<@O             `@
                           �?9'���l	@�           4�@                          �:@�^���		@Q            @`@������������������������       �*�/}�&@@            @Y@������������������������       ��sᜨ�@             =@                            �?Jq���H	@�           ,�@������������������������       ��1�*�@           �z@������������������������       �Uh_�@r	@           ��@                           @�s���@J           P�@                           @�U���@           p�@                           @1j�x�@            z@������������������������       �֯���O@�            �r@������������������������       �(6x0�@@            @]@                            �?O���� @�           ��@������������������������       ��S�-sa @           �{@������������������������       �G��{�9@�            x@                            �?�����@E           �@                           �?�$S6�@P             `@������������������������       ���}�j@(            @P@������������������������       ��ΙOdI@(            �O@                          �5@�ȑ�2V@�            �w@������������������������       ���ۘ��@�            `k@������������������������       ���CE'�@e            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �s@     `�@      >@     �N@     �|@     @T@     ��@     �j@      �@     �s@      <@      6@     �l@     �s@      8@     �D@      t@     �P@     �v@     �e@      w@     @k@      3@      �?      R@      R@      �?      $@     @R@      @     `f@      ;@     @_@      H@      @      �?      .@      6@              @      0@       @     �N@      @     �H@      "@       @      �?      @      &@              @      &@       @      @@      @      .@      @                      &@      &@                      @              =@       @      A@       @       @             �L@      I@      �?      @     �L@      @     �]@      6@      S@     �C@      �?             �B@     �E@      �?      @     �E@       @     �Q@      2@      G@      A@      �?              4@      @                      ,@      �?      H@      @      >@      @              5@     �c@      n@      7@      ?@      o@     �N@     �g@     �b@     �n@     @e@      0@      @      *@      2@              @      9@      @      @      8@      0@      *@      @      �?      "@      *@              @      9@      �?      @      3@      .@      "@               @      @      @                               @              @      �?      @      @      2@      b@     �k@      7@      :@      l@      M@      g@      _@     �l@     �c@      $@      @      G@     �P@      @      @     @P@      1@     �Q@     �J@      P@      A@       @      .@     �X@     �c@      4@      6@     �c@     �D@     @\@     �Q@     �d@     �^@       @       @      U@     �j@      @      4@     �`@      .@     Ѕ@      C@     �z@     �X@      "@       @      K@     �b@      �?      @      V@      &@     ��@      4@     0s@     �N@      @       @      7@      L@      �?      �?      @@      &@     �c@      *@     �U@      @@      @       @      $@      D@              �?      7@      "@     @`@      @      M@      5@                      *@      0@      �?              "@       @      :@       @      <@      &@      @              ?@      W@              @      L@              x@      @     �k@      =@       @              (@      H@                      A@             @i@      @     �_@      ,@                      3@      F@              @      6@             �f@      �?     �W@      .@       @              >@      P@      @      *@     �G@      @     �c@      2@     �^@      C@      @               @      @              �?       @      @     �H@      @      D@      $@                      @      �?              �?      @      �?      5@       @      5@       @                      @      @                      @       @      <@      �?      3@       @                      6@      M@      @      (@     �C@      �?     @[@      .@     �T@      <@      @              1@     �C@       @      @      ,@      �?      T@      @      F@      @      @              @      3@      @      @      9@              =@      $@     �C@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�J6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@X�#>�*@�	           ��@       	                    @���n�q@�           l�@                          �0@�q�^�@-           }@                           @2ħve@4             S@������������������������       ��w�~h@'             L@������������������������       ��Dá� @             4@                          �1@E�)7��@�            Px@������������������������       �r���d@u            �g@������������������������       ���b�:�@�             i@
                           @u_�1�H @T           P�@                           @���-r�?           @|@������������������������       ��<%Q���?�            �m@������������������������       ���ɝ�� @{             k@                           �?� �s&@@Q            �`@������������������������       ��	���?(            �P@������������������������       ��ƃ��s@)            �P@                            @$�o��@0           \�@                          �7@w��p�@            �@                          �5@M��{F�@%           ��@������������������������       ��l4L�5@6           h�@������������������������       �}��$��@�            @w@                          �:@�<�H�@�           ��@������������������������       ����;�@�             x@������������������������       ��V��Xa@�            �y@                           @���D�@           p�@                          �<@܉�s�L	@�            �@������������������������       ����Κ�@Z           h�@������������������������       ��[�)U�	@F            �\@                           �?S���@u            �e@������������������������       �I�W@7            �T@������������������������       ���eg�@>            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     q@     Ё@     �C@      G@     �~@      T@     ��@     �i@     �@      u@     �@@      �?      E@     @`@              @     �Y@       @      {@      B@     �j@     �T@      �?      �?      7@      P@              @     �Q@      @     �`@      >@     @T@     �K@      �?              @      3@               @      .@              2@      @       @      @                       @      &@               @      ,@              *@       @       @      @                      @       @                      �?              @      @                              �?      2@     �F@              �?     �K@      @     �\@      9@     @R@     �I@      �?               @      6@                      3@      �?      P@      *@     �D@      4@              �?      $@      7@              �?      B@      @      I@      (@      @@      ?@      �?              3@     �P@                      @@      @     �r@      @     �`@      ;@                      0@      I@                      &@      @      o@      @      Y@      4@                       @      >@                      �?      @     �b@      �?      D@      @                       @      4@                      $@             �X@       @      N@      1@                      @      0@                      5@             �I@      @     �@@      @                              *@                       @             �@@              *@                              @      @                      *@              2@      @      4@      @              0@     �l@     �{@     �C@     �E@      x@      R@     ��@     `e@     8�@      p@      @@       @     �c@     0s@      5@      =@     pq@     �N@     �}@      \@     py@     �e@      5@      @     @V@      i@      ,@      0@     �c@      =@     �u@     �K@     0p@     @Q@      "@      @     �F@     �b@      @      $@     @Z@      4@     `o@      C@      h@     �J@      @      �?      F@     �I@       @      @     �J@      "@     �W@      1@     �P@      0@      @      @     �Q@     �Z@      @      *@     @^@      @@     �_@     �L@     �b@     �Y@      (@             �B@      P@       @      &@     �F@      0@     @P@      4@      S@     �C@      "@      @     �@@     �E@      @       @      S@      0@     �N@     �B@      R@      P@      @       @      R@     �`@      2@      ,@     �Z@      &@      c@     �M@      b@      U@      &@       @     @Q@     �]@      2@      ,@     �V@      "@     @T@     �L@     �W@      R@      "@      @      K@     �Y@      *@      @     @R@      @     @S@     �D@     �U@      K@      "@      @      .@      1@      @       @      1@      @      @      0@       @      2@                      @      ,@                      1@       @      R@       @      I@      (@       @              �?      "@                      @              A@      �?      :@      @       @               @      @                      &@       @      C@      �?      8@       @        �t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�K\bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�,Wf�+@�	           ��@       	                   �<@կc�@           �@                           �?NGrHy�@�           ��@                           �?�+����@           �y@������������������������       �2��z@i            �d@������������������������       �k
%��@�            �n@                            �?�2�}}@�           X�@������������������������       �ϒn�<j�?w            �f@������������������������       ��:YHQl@W           ��@
                           @�~���@=            �X@                           �?����X�@2            @T@������������������������       �I��~!�@             D@������������������������       �CtmR�&@            �D@������������������������       �ѥA��@             2@                           @;�A4	@�           �@                           @��H}�	@�           ��@                           �?}1!kKU	@l           p�@������������������������       ����$��@L            @^@������������������������       �!�S�;3	@            ��@                           �?$����Y	@Y           ��@������������������������       ��
�	@�            x@������������������������       �"-��@\            �c@                          �7@O*��d@�           X�@                           @�X
9	C@"           0�@������������������������       �;߼�z@           Ȋ@������������������������       �YL��J@             *@                           @���dj@�             s@������������������������       � ��B.@�             o@������������������������       �5�5��;@             L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     `r@     ��@      <@     �M@     �|@     �Q@     H�@      j@     Ј@      w@      @@              X@     �f@              &@     �X@      &@     �z@      A@     Pq@      U@      @             �T@     �d@               @     �U@      $@     �y@      =@     �p@      M@      @              H@      R@              @     �J@      @     �W@      6@     @T@      :@      @              @      >@                      3@              L@      @      C@      @      �?             �D@      E@              @      A@      @      C@      0@     �E@      3@       @             �A@      W@              @     �@@      @      t@      @     `g@      @@      �?              �?      .@              �?      @              Y@              J@      @                      A@     @S@               @      :@      @     �k@      @     �`@      :@      �?              *@      0@              @      *@      �?      *@      @      "@      :@                      *@      (@              @      (@              @      @       @      9@                      @       @               @       @               @      @       @      1@                      "@      @              �?      $@               @      �?      @       @                              @                      �?      �?      "@      �?      �?      �?              0@     �h@     @v@      <@      H@     �v@      N@     8�@     �e@     (�@     �q@      <@      0@     ``@     �j@      9@     �D@     0p@     �F@      j@      b@     `k@     `g@      9@      ,@     @W@     �]@      .@      8@     �f@      ?@      `@     @Q@     `c@     ``@      *@      @      $@       @              @      <@       @      @      (@      3@      5@      @      "@     �T@     �[@      .@      2@     @c@      =@     @^@     �L@      a@     �[@      $@       @      C@      X@      $@      1@     @S@      ,@      T@      S@      P@      L@      (@       @      ?@     �L@      @      ,@     �L@      $@     �I@      N@     �B@     �G@      (@              @     �C@      @      @      4@      @      =@      0@      ;@      "@                     �P@     �a@      @      @      Z@      .@     py@      >@     �r@     �X@      @              H@     �\@              @      N@      *@     �t@      *@     @l@     �N@      �?              G@     �\@              @     �M@      $@     `t@      *@      l@     �M@      �?               @                              �?      @      @              �?       @                      3@      :@      @      @      F@       @     @S@      1@      R@      C@       @              $@      5@      �?      @      D@              Q@      (@      M@      A@                      "@      @       @              @       @      "@      @      ,@      @       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��LhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�&/ȟ@�	           ��@       	                    �?'��>u	@�           ��@                          �<@��@*��@           �x@                           �?�ϮEՆ@�            �u@������������������������       �O+1��@l            `b@������������������������       �7B�-@�            �h@                           �?AuN��@#            �J@������������������������       ��d�1� @
             .@������������������������       �F:8`��@             C@
                           �?�>���	@�           \�@                          �3@����&@            {@������������������������       � �:���@Y             b@������������������������       �Z���.@�            �q@                          �;@f�}�S
@�           8�@������������������������       ����	@j           x�@������������������������       ��m��	@[             c@                          �5@h)����@�           F�@                           @���@�           x�@                           @�9^'@�            �u@������������������������       �+��+��@X             b@������������������������       �W�
���@            �i@                          �4@�(7��@�           �@������������������������       ��,=e@T           �@������������������������       �QgQPZ�@b            �c@                          �=@m�ckQ�@%           (�@                           �?��̙4@�           P�@������������������������       ��_%)�m@�            �i@������������������������       ���֢0�@p           ��@                           @DxF9�f@5            �V@������������������������       �8��@#            �M@������������������������       ��8�Rj@             @@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@      u@     ��@      @@     �L@     �}@      U@      �@     �l@     ��@     0u@     �D@      2@     �e@     �m@      7@     �@@     @p@      H@      j@     �_@     @n@     �e@      @@       @      F@     @Q@      �?      @     �J@      @     �S@      4@      T@      F@      �?       @      E@      L@      �?      �?     �E@      @      S@      1@     @S@      :@      �?       @      0@      5@      �?      �?      3@      @      ?@      $@      >@      (@                      :@     �A@                      8@             �F@      @     �G@      ,@      �?               @      *@               @      $@               @      @      @      2@                       @      @                       @              �?                      @                              @               @       @              �?      @      @      .@              0@     @`@     �d@      6@      >@     �i@      F@     ``@     �Z@     @d@      `@      ?@              7@      O@      @      *@     @U@       @     �S@     �F@      O@      G@      @              .@      1@                      3@      �?     �A@      2@      8@      .@      �?               @     �F@      @      *@     �P@      @      F@      ;@      C@      ?@      @      0@     �Z@     @Z@      1@      1@     �^@      B@      J@     �N@      Y@     �T@      ;@       @     �S@     �R@      "@      (@     @[@      5@     �I@     �J@     @U@     �P@      8@       @      =@      >@       @      @      *@      .@      �?       @      .@      1@      @      @     @d@     0u@      "@      8@      k@      B@     ��@     �Y@     P~@     �d@      "@             �I@      k@      @      *@      \@      $@     (�@      H@     �s@      T@      @              .@      Q@      �?      @     �A@      @     �\@      B@     �K@      .@                       @      &@               @      4@      �?      O@       @      7@      "@                      @     �L@      �?       @      .@      @     �J@      <@      @@      @                      B@     �b@      @      "@     @S@      @      }@      (@     @p@     @P@      @             �@@     @^@      @       @     �K@      @     @z@      &@     �j@      O@      �?              @      <@              �?      6@      @      G@      �?      G@      @      @      @     �[@     �^@      @      &@     @Z@      :@     �i@      K@     @e@     �U@       @      @     �V@     �Z@      @      "@      W@      2@     `h@      I@     �d@     @S@      �?              $@      4@      �?              &@      @     �U@       @     �K@      ,@              @     @T@     �U@      @      "@     @T@      *@     @[@      H@     @[@     �O@      �?              4@      0@      �?       @      *@       @      &@      @      @      "@      �?              ,@      @               @       @      @      "@      @       @      "@      �?              @      $@      �?              @      @       @              @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ �hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?8�#B"C@�	           ��@       	                    �?w�&{&@            �@                           �?�ń\)@~           ��@                           �?�7�'a@�            @k@������������������������       ��ٙ��S@8            �U@������������������������       ��Bz�:�@S            �`@                          �:@���~� @�            @x@������������������������       ���C6�I @�            @u@������������������������       ��h��dA@             H@
                          �<@�_��7@�           P�@                           �?{1_�l@g           �@������������������������       �I=p�<@�            �m@������������������������       ���$F�a@�            u@                          �@@���o@             �F@������������������������       ��6�k�@             B@������������������������       �R�F V�?             "@                          �5@nc!KC@�           �@                           @�a	U5�@~           �@                           @����q�@E           ��@������������������������       ��;A~F@"            ~@������������������������       �D�K@#            }@                           �?<k��\@9           @�@������������������������       �m����@�            `l@������������������������       ��e�NI@�            Pr@                          �<@�ƾ��V	@           �@                           �?��}��	@t           ��@������������������������       ����d@�            @y@������������������������       �].?��b	@w           �@                           �?y��!G	@�            �m@������������������������       �v��RA�@             9@������������������������       ��d�.	@�            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@     �@@     �G@     `{@      R@     ��@     p@     ��@     �t@      A@       @      T@     @f@       @      @     @W@      "@     �{@      F@     �r@     �Q@       @       @     �A@      S@       @      @      E@      @     �m@      2@     �a@      E@               @      :@      B@       @      @      4@       @     �E@      *@      H@      6@               @      @      @                      &@              8@      @      ;@      @                      5@      =@       @      @      "@       @      3@      $@      5@      .@                      "@      D@               @      6@      @     @h@      @      W@      4@                      @      ?@               @      6@      @      f@      @      T@      ,@                       @      "@                              �?      1@      �?      (@      @                     �F@     �Y@              �?     �I@      @     �i@      :@     �c@      <@       @              D@      X@                      E@      @      i@      7@     �b@      3@       @              7@      D@                      =@              N@      .@     �K@      (@       @              1@      L@                      *@      @     �a@       @     @W@      @                      @      @              �?      "@              @      @       @      "@                      @      @                      @              @       @       @       @                              �?              �?      @                      �?              �?              0@      m@     �u@      ?@      D@     �u@     �O@     (�@     �j@     x�@     0p@      @@      @     �V@      i@      $@      3@      f@      ?@     �x@     �U@     �t@     �\@      *@       @     �K@     �^@      @      $@     ``@      9@     �n@     �M@     �k@     @Q@      �?       @      B@      N@      @      "@     �U@      1@     �V@      H@     �T@     �F@      �?              3@      O@      �?      �?     �F@       @     `c@      &@     �a@      8@               @      B@     �S@      @      "@     �F@      @     �b@      <@     @Z@     �F@      (@      �?      1@     �E@      @      @      3@      @     �N@      (@     �A@      4@      @      �?      3@      B@              @      :@       @      V@      0@     �Q@      9@      @      (@     �a@     �b@      5@      5@      e@      @@     `g@     �_@     �h@      b@      3@      $@      \@     �\@      ,@      0@      a@      4@     @e@     @W@     `e@     �Z@      3@              E@      M@      @       @     �L@       @      P@      @@     �R@     �K@      &@      $@     �Q@      L@      @      ,@     �S@      2@     �Z@     �N@     @X@      J@       @       @      =@     �A@      @      @     �@@      (@      1@     �@@      <@      C@                      @      @              @      @                      @      �?       @               @      :@      =@      @       @      =@      (@      1@      ;@      ;@      B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ2&hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�f���m@�	           ��@       	                   �3@��&y�@p           8�@                            �?��T�@�           �@                          �0@	�O�J�@�            �l@������������������������       �5��\��@             E@������������������������       ����kn@o            �g@                           �?1���@B           �@������������������������       �8�rnm�@s            @f@������������������������       ��E��l@�            �t@
                           �?�-L��`	@�           �@                           �?d,f夅	@�           ��@������������������������       �o�k��@�            s@������������������������       �/�D�Y�	@           �@                           �?[z�V�K@�            �t@������������������������       �b��Y��@6            �T@������������������������       ��_v�M�@�            @o@                            @�Hw�^@:           ��@                           @������@�           P�@                           @����q@}           ؎@������������������������       �1��Ov@�            �t@������������������������       ��{����@�           ��@                            �?�1��@           �{@������������������������       ��T�ݟ+@�            Pt@������������������������       ��m|>xy@I             ]@                           @�oh�>�@�            �q@                           @��,�w% @\            `b@������������������������       �ؒ�NW @O            �_@������������������������       �:�~t��?             5@                           �?Z#����@U            �`@������������������������       ��\�#
@)             O@������������������������       �q�񡃼@,             R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      r@     ��@      ;@     �K@     �|@     �V@     ��@     `l@     @�@     v@      >@      7@     @j@     �u@      6@     �C@     �t@     �N@     x@     `f@     �u@     �m@      9@      @     �G@     @Y@      @      @     @W@      &@     �h@     �M@     �b@     �N@      @              ,@      ?@                      :@      �?     �O@      4@      O@      ,@                      @      "@                      @              1@      �?       @       @                       @      6@                      5@      �?      G@      3@      N@      (@              @     �@@     �Q@      @      @     �P@      $@     �`@     �C@      V@     �G@      @              3@      <@                      4@       @     �K@      @      D@      @              @      ,@      E@      @      @     �G@       @     �S@      @@      H@      D@      @      1@     `d@     �n@      0@     �A@     `m@      I@     �g@      ^@      i@     �e@      6@      1@     @]@     �g@      ,@      9@     `h@      D@     �`@     �W@     �a@     �a@      5@      �?      @@     �L@      @      "@      B@       @     �L@      8@      J@      >@      �?      0@     @U@     �`@      $@      0@     �c@      C@     �S@     �Q@     �V@     @\@      4@              G@     �J@       @      $@      D@      $@      K@      :@     �M@      @@      �?              ,@      @                      (@              >@      @      *@      @                      @@     �G@       @      $@      <@      $@      8@      7@      G@      ;@      �?      �?      T@     �k@      @      0@     �`@      >@     ��@      H@     �|@     @]@      @      �?     �Q@     `i@      @      &@     �[@      =@     ~@      F@     Pw@     @X@      @      �?      E@     �a@              @     �Q@      1@     �v@      5@      p@     �P@      �?      �?      .@     �K@              �?      9@      0@     �Z@      $@     �P@     �@@      �?              ;@     �U@               @     �F@      �?     @p@      &@      h@      A@                      =@      O@      @       @      D@      (@     �\@      7@     �\@      >@       @              5@     �D@      @      @      A@      $@     @V@      $@      U@      :@                       @      5@       @      �?      @       @      :@      *@      ?@      @       @              "@      4@              @      7@      �?     @\@      @      U@      4@       @               @      $@                      .@             �M@      �?      K@      @       @              �?      "@                      .@              L@      �?      C@      @       @              �?      �?                                      @              0@                              @      $@              @       @      �?      K@      @      >@      0@                       @      @               @      @      �?      9@              *@      $@                      @      @              @      @              =@      @      1@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ"�YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��7f�M@�	           ��@       	                    �?����?�@x           $�@                          �7@>�K'@�           ��@                           �?�Y��e@           �x@������������������������       ��j���@|            @g@������������������������       �2T����@�            �j@                            @��0�� @�            @m@������������������������       �k߫�_�@Z             b@������������������������       ��ƺG�@5            @V@
                          �3@R��у	@�           h�@                           �?��I1'@(           P}@������������������������       ��'�:��@�            ps@������������������������       ��s��Z�@c            �c@                           �?"A���	@�           �@������������������������       ���V@�            pq@������������������������       �?�+��	@           p�@                            @}ўQ��@F           ܚ@                            �?���@�           ��@                           @�>���@j           ��@������������������������       ���P\��@_           �@������������������������       ���˓�@             .@                          �4@���|u@;           0@������������������������       ���M�L@�            0q@������������������������       �]ɗ�Ɇ@�             l@                           @�8ha]@�             q@                          �3@����'�?\            �c@������������������������       �D��J���?,            �Q@������������������������       ���(	�?0            �U@                           @���yR�@E            @]@������������������������       �r _��}@8            �W@������������������������       ��� A�@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      s@     @�@      A@     �M@     �|@     �V@     �@     �l@     h�@      u@      8@      .@     �j@     �r@      9@     �G@     �t@      Q@     pw@     �f@     �w@     `l@      8@       @      L@     �R@       @      $@     �U@      @      e@      @@     `c@      D@      @             �B@      F@              @      D@      �?     �_@      0@     �Z@      5@                      &@      :@              @      4@      �?      Q@      $@      B@      $@                      :@      2@              �?      4@             �M@      @     �Q@      &@               @      3@      >@       @      @      G@      @     �D@      0@      H@      3@      @       @      ,@      3@              �?      6@      @      =@      @      >@      0@      @              @      &@       @      @      8@              (@      $@      2@      @              *@     �c@     �l@      7@     �B@     �n@      P@     �i@     �b@     �l@     `g@      5@      @     �A@     �O@      @      @      P@      "@     �Y@     �E@     �R@     �M@      @      @      >@     �D@      @      @      E@      @      K@      ?@      H@     �E@      @              @      6@              @      6@       @     �H@      (@      ;@      0@              $@      _@     �d@      2@      >@     �f@     �K@      Z@     @Z@      c@      `@      2@              9@     �H@       @      $@     �I@      @     �C@      ,@      E@     �B@      @      $@     �X@      ]@      0@      4@     �`@     �I@     @P@     �V@     �[@     �V@      (@      @     @V@     @k@      "@      (@     @_@      6@     p�@      H@     �z@     @[@              @     @S@     �h@      @      "@     @[@      2@     x�@      F@     �v@     �W@                     �D@     @_@       @      @      T@      (@     �u@      ;@      n@     @P@                      C@     @_@      �?      @     �S@      "@     �u@      ;@     �m@     @P@                      @              �?       @      �?      @      �?              @                      @      B@     @R@      @      @      =@      @     �f@      1@      ^@      =@                      &@      E@              @      @      @     �`@       @     �N@      "@              @      9@      ?@      @              7@      @      H@      "@     �M@      4@                      (@      4@      @      @      0@      @     �_@      @     @Q@      .@                       @      &@                      $@             �S@      �?      G@       @                       @      &@                      @             �@@      �?      5@                              @                              @              G@              9@       @                      @      "@      @      @      @      @      H@      @      7@      *@                      @      @              @      @              E@      @      5@      (@                              @      @               @      @      @               @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�X�vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @"u��v@�	           ��@       	                    �?#�D�		@~           ��@                            �?͚�yNi	@	           Й@                           �?�?�w}�@B           �@������������������������       ��s��s@f            �c@������������������������       ���B	@�            �u@                           �?��Z��	@�           �@������������������������       ��E���	@            z@������������������������       ��t w=7	@�           І@
                          �4@�G
=�K@u           ��@                            �?Y�.a��@�            0r@������������������������       ��G	{@l             g@������������������������       �}�r�e@E            �Z@                           �?���X@�             s@������������������������       ��T;��@2            @R@������������������������       ��k�S'�@�            �l@                          �5@���|��@<           �@                          �1@��ʷo@�           �@                           @AxG߇��?�            �s@������������������������       �&Ek���?�            �o@������������������������       ��J��k@-            �P@                           �?�o��`O@�           8�@������������������������       � m����@�            @w@������������������������       �?0}��/@�            0u@                            @���섬@�           ��@                          �6@�Mw>�@R           h�@������������������������       ����̚s@;            @W@������������������������       ���2)@            {@                           �?gN���@D            �[@������������������������       ��B�M� @             H@������������������������       ��;�F2� @%            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @s@     Ѐ@      A@     �M@     `|@     �W@     �@     `i@     `�@     �v@      ?@      5@     �k@     `s@      <@     �E@     �t@     @R@     �w@     `e@     @x@     0p@      ;@      5@     �d@     �k@      ;@     �B@      o@      H@     �n@      _@     �p@      k@      :@      "@     �K@     @Q@      �?       @     @T@      "@     �U@      F@     @V@      F@      $@       @      .@     �A@              �?      1@              C@      @     �A@      @       @      @      D@      A@      �?      @      P@      "@      H@      D@      K@     �B@       @      (@     �[@      c@      :@      =@      e@     �C@     �c@      T@     �f@     �e@      0@      @      F@      O@      0@       @     �L@      4@      L@      6@      J@     @Q@      @      @     �P@     �V@      $@      5@     �[@      3@     �Y@      M@     @`@     �Y@      &@              L@      V@      �?      @     �S@      9@     �`@     �G@     @]@     �E@      �?              ,@     �G@      �?              C@       @     @T@      1@     @Q@      6@                      (@      :@      �?              4@       @     �K@      (@     �C@      1@                       @      5@                      2@              :@      @      >@      @                      E@     �D@              @     �D@      7@     �I@      >@      H@      5@      �?              @      $@                      "@      @      7@      @      ,@      �?      �?             �A@      ?@              @      @@      2@      <@      ;@      A@      4@                     �U@     �l@      @      0@     �_@      6@     @�@      @@     �z@     �Z@      @              C@     `a@      @      &@     �Q@       @     �z@      "@     0q@      G@      @              @      D@              @      1@             �c@      �?     @T@      &@      �?              @      =@                      "@              a@             �P@      @                      �?      &@              @       @              7@      �?      ,@      @      �?             �@@     �X@      @      @     �J@       @     �p@       @     @h@     �A@       @              *@      H@      @      @      F@      @      a@      @      W@      6@      �?              4@     �I@              @      "@      @     ``@      @     �Y@      *@      �?              H@     @V@       @      @      L@      ,@     �g@      7@     �b@      N@      �?             �E@     �T@      �?      @     �H@      ,@     �b@      7@     �[@      I@      �?               @      &@      �?              "@      @     �D@               @      (@                     �A@     �Q@              @      D@      &@      [@      7@     �Y@      C@      �?              @      @      �?       @      @              D@             �C@      $@                              @               @       @              3@              .@      @                      @              �?              @              5@              8@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?R�S�L-@�	           ��@       	                    �?���jļ@           ��@                           �?t>V��@�           �@                            �?�񣷡^@�            @j@������������������������       �2�rt��@&             O@������������������������       �~V��o@d            �b@                           @�`&��(@           {@������������������������       ��z��U;@�             s@������������������������       �>W1Wݫ@N            �_@
                          �5@�i�u�G@t           X�@                            �?�C��dB@�             x@������������������������       �0zY�ڟ�?<             Y@������������������������       �rRE, j@�            �q@                          �<@��CT@�            `m@������������������������       ��Va��@o            @f@������������������������       ��|�h�@"            �L@                           �?�V�
@�           ��@                           �?�,��	@�           X�@                           �?� �׍�@�            �x@������������������������       �[�E�R!@]            @a@������������������������       �*M��E@�            0p@                            @�[!z�	@�           H�@������������������������       �3-D^�n
@           �y@������������������������       ��C�W�@�            s@                          �6@x�\���@�           �@                           @ 4�1p�@�           ��@������������������������       �吺P4�@�            @r@������������������������       ����J�@�           `�@                            �?���8@K           ��@������������������������       ��."�
@]            �b@������������������������       �����`@�            �w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �q@     0�@      6@      P@     �{@      U@     ��@     `m@     `�@     �s@      8@      �?     �R@     �c@       @      (@     �]@      1@     �{@     �L@     ps@     �P@      @      �?      D@      Q@       @      &@      J@      *@     @o@      A@     �a@      >@       @      �?      .@      <@       @      @      :@      @      G@      7@      D@      .@       @      �?      �?      @              @      &@      �?      .@      "@      &@      @                      ,@      5@       @      @      .@      @      ?@      ,@      =@      (@       @              9@      D@              @      :@       @     �i@      &@      Y@      .@                      2@      >@              �?      0@      @     �b@      "@     �Q@      @                      @      $@              @      $@      @     �J@       @      =@      $@                      A@      V@              �?     �P@      @      h@      7@     `e@      B@      @              1@      G@              �?      =@              c@      @     �[@      4@       @              �?      .@                                      J@              >@       @                      0@      ?@              �?      =@              Y@      @      T@      2@       @              1@      E@                     �B@      @      D@      0@     �N@      0@       @              &@     �A@                      9@      @     �A@      @     �J@       @      �?              @      @                      (@              @      $@       @       @      �?      8@     �i@     �x@      4@      J@     �t@     �P@     (�@     @f@     ��@     @o@      2@      7@     @\@     `e@      (@      :@     `f@      D@      `@     @\@     �d@     �^@      1@      @      7@     @Q@      �?      $@     �N@      "@      R@     �A@      P@      E@      @      @      "@      9@              @      A@      @      4@      *@      ,@      (@       @      @      ,@      F@      �?      @      ;@      @      J@      6@      I@      >@      @      1@     �V@     �Y@      &@      0@     �]@      ?@     �L@     �S@      Y@     @T@      (@      "@     �K@      H@      @      &@     �M@      6@     �@@      J@     �G@      K@      &@       @     �A@      K@      @      @     �M@      "@      8@      :@     �J@      ;@      �?      �?     @W@     �k@       @      :@     �b@      ;@     @|@     @P@     w@     �_@      �?              J@      b@      @      1@      T@      0@     �u@      >@     �n@      R@                      $@      H@       @      &@      ?@      @     @T@      7@     �M@      6@                      E@      X@      @      @     �H@      &@     �p@      @      g@      I@              �?     �D@     �S@       @      "@     @Q@      &@     @Z@     �A@     @_@     �K@      �?              (@      6@               @      ,@      @      F@      @      @@      0@      �?      �?      =@     �L@       @      @     �K@       @     �N@      >@     @W@     �C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJWV�RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�`1�$e@�	           ��@       	                    �?�,�O�@k           ,�@                           �?�ty%^@�           �@                          �<@��	I�@H           �@������������������������       ��zq@            �{@������������������������       �S���Z�@(             N@                            �?�
n�A�@y             i@������������������������       ���<E�@.            @R@������������������������       �Y�YP�@K            �_@
                           �?~�7�Mr	@�           P�@                           �?�a���	@�           0�@������������������������       �~���K�@           �z@������������������������       ��\z�O
@�           �@                          �1@�Z�IS�@�            �x@������������������������       ��K:�d@%            @P@������������������������       �����K@�            pt@                          �4@m��`ta@2           ̚@                           �?p�S#�@9           ؋@                            @p�]Ʋ�?�            �t@������������������������       �=�AQ�S�?�            `p@������������������������       ����8<�?'             Q@                           @h^��/�@f           ��@������������������������       ����"?@=            �V@������������������������       ��{�F1@)           p}@                           @��
�Rs@�           ��@                           @�-�*��@G            �@������������������������       �\w���q@            `~@������������������������       �13E�{@'             M@                            @�	V�)z@�            �q@������������������������       ����Z@�            �l@������������������������       �nN���@$             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     ��@     �A@     �J@     `{@      S@     P�@      m@     ��@      x@     �@@      2@     �j@      t@      7@     �C@     �r@     �K@     px@     @g@     �v@     �p@      ;@      �?      R@     �W@      @      "@      S@      @      g@      B@     �d@     �L@      @      �?     �I@     �S@      @      @      P@       @     @]@      ;@     �Y@     �H@      @      �?      F@     @Q@      @       @      L@       @     �\@      8@     �W@      ?@      @              @      $@              @       @              @      @       @      2@                      5@      .@              @      (@      �?      Q@      "@     �N@       @      �?              @       @              @      @      �?      5@              9@       @      �?              0@      @                      @             �G@      "@      B@      @              1@     �a@     �l@      4@      >@     �k@      J@     �i@     �b@     �h@      j@      5@      1@     @^@     �b@      4@      :@      e@     �E@      `@     @Z@     @a@      d@      5@              ?@      M@      @      ,@     �O@      (@     @S@     �A@      L@     �P@      @      1@     �V@     @W@      ,@      (@     �Z@      ?@     �I@     �Q@     �T@     �W@      ,@              6@     @S@              @     �I@      "@     �S@     �F@     �M@     �G@                              ,@                      @              8@      (@      @      @                      6@     �O@              @     �G@      "@      K@     �@@      J@     �E@              @     @P@     �n@      (@      ,@     �a@      5@     �@      G@     �z@     @^@      @              <@      ^@      @       @      B@       @     @y@      ,@     @l@     �H@                      "@     �B@              �?      "@             �g@      �?     @R@      &@                      @     �B@                       @              b@      �?     �K@      $@                      @                      �?      �?              F@              2@      �?                      3@     �T@      @      @      ;@       @     �j@      *@      c@      C@                      @      2@              @      @              7@      @      6@      "@                      .@     @P@      @      �?      7@       @      h@      "@     ``@      =@              @     �B@     �_@       @      @     �Z@      3@     �i@      @@     @i@      R@      @      @      6@     �S@      �?       @     �Q@      "@     �c@      .@     �`@      G@      @      @      1@     �P@               @      N@      @     `b@       @     �`@      E@      �?              @      &@      �?              &@       @      "@      @      @      @      @              .@      H@      @      @     �A@      $@     �I@      1@     �P@      :@                      ,@     �D@      @       @     �@@      $@      B@      ,@      L@      1@                      �?      @       @       @       @              .@      @      &@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�/gchG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���[A@�	           ��@       	                   �<@㭋K�@           В@                           �?�vF �3@�           |�@                           �?M�^��@�             y@������������������������       ��9�T�-@s             h@������������������������       �H���@�            �i@                            �?��$��@�           x�@������������������������       ��>�9Pr�?o            �d@������������������������       ���3x�j@]           H�@
                           �?TL�� @9            @U@                           �?9�Vw�@            �H@������������������������       �>��_�@
             0@������������������������       �ϻ���@            �@@                            �?�>zA�E@             B@������������������������       �hJN�@             "@������������������������       �.�)�,@             ;@                           @h��zk@�           *�@                           �?eF�j9	@�           ԗ@                           �?���s�{	@�           ,�@������������������������       �4dr�|@           �y@������������������������       �\�8�	@�           `�@                          �4@��s@           �z@������������������������       ����R�@p            �e@������������������������       ��R���@�            �o@                           @�Hx�@�           ��@                          �<@�R�65@}           0�@������������������������       �m1���@X           ��@������������������������       �����v@%             L@                            �?��|I@X            �b@������������������������       �q�ړ@             I@������������������������       �t�m��@@            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     p�@      <@     �F@     p~@     �R@     p�@     `l@      �@     �u@     �@@       @      T@     �c@       @       @      ]@      (@     `z@     �D@     0q@     �S@      @       @      S@     @b@       @      �?     �Z@      &@     �y@      ?@     �p@      O@       @       @     �D@     �M@       @             �I@      @     @W@      7@     �T@     �B@      �?       @      6@      2@       @              :@      @     �K@      &@      @@      0@                      3@     �D@                      9@              C@      (@      I@      5@      �?             �A@     �U@              �?     �K@       @     �s@       @      g@      9@      �?                      5@              �?      "@      �?     @V@             �C@      @                     �A@     �P@                      G@      @     @l@       @      b@      3@      �?              @      (@              @      $@      �?      ,@      $@      "@      1@      �?              @      @              @       @              @      @      @      (@                       @      @                      �?              @               @      @                       @      @              @      @                      @      �?       @                              @                       @      �?      &@      @      @      @      �?                      �?                       @      �?               @       @              �?                      @                                      &@      @      @      @              *@     �m@      y@      4@     �B@     0w@      O@     @�@     @g@     @      q@      >@      *@     �c@     �l@      (@      >@      o@     �K@     �k@     @c@     �i@     @f@      7@      *@      _@     @c@      $@      7@     �g@     �B@      a@     �[@     `b@     �`@      6@      �?      9@     �P@       @      ,@     �R@      @     �P@      D@     �M@     �J@      @      (@     �X@      V@       @      "@     �\@      >@     @Q@     �Q@      V@     @T@      .@             �A@     �R@       @      @     �N@      2@      U@     �E@     �L@      F@      �?              @      E@       @              1@      �?     �J@      ,@      7@      1@                      @@      @@              @      F@      1@      ?@      =@      A@      ;@      �?             �S@     �e@       @      @     �^@      @     �v@      @@     Pr@     �W@      @              N@     �b@      @      @      \@      @     �t@      8@     �p@     �Q@                     �J@     �a@      @      @     �W@      @     �t@      8@     `p@     �N@                      @       @              �?      1@              @               @      $@                      2@      8@      �?       @      $@      @      =@       @      7@      7@      @              @      @      �?       @                       @       @      "@      .@                      &@      2@                      $@      @      5@      @      ,@       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@+��B�X@�	           ��@       	                   �1@\����@C           ��@                           �?�X�xG�@�           ��@                           �?sf�L�@l            �e@������������������������       �d�ݫ��@1             T@������������������������       ��9� ��@;            �W@                           @Z���q@           `|@������������������������       ��ߍ���?�            �v@������������������������       ��[��_i@6            �W@
                           @ً6"��@�           ��@                           �?����
@           ؉@������������������������       �u�:��P@i           ��@������������������������       �bdϩ�@�            �l@                           @���%�N@�           h�@������������������������       �")ܴ�q@8           �~@������������������������       �Xu����@�            `h@                           �?�՞�X�@N           ��@                            �?י^�Zi@           }@                           �?���3��@Q             ^@������������������������       ���cc @5            �T@������������������������       ��d�(�@             C@                           �?�0|2��@�            �u@������������������������       �9����X@n            @f@������������������������       ��v��@_            �d@                          �:@�Ro�	@0           l�@                          �9@���5�]@           �@������������������������       �q��3�@�           p�@������������������������       �=�ա�X@X            �a@                            @����M	@           �{@������������������������       ��=�4P@�            �q@������������������������       �FM��Y�	@\            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �t@     ��@      2@      K@     �|@      T@     ��@      l@     8�@     �w@      ?@      @     �a@     �s@      @      =@      g@      ;@     0�@     �W@     �|@     �g@      &@      �?      ?@      S@      �?      $@     �D@             �o@      5@     �b@      F@       @      �?      1@      4@      �?      @      5@              C@       @     �C@      :@              �?      @      "@      �?               @              4@      @      (@      4@                      *@      &@              @      *@              2@      @      ;@      @                      ,@      L@              @      4@             �j@      *@     �[@      2@       @               @     �C@                      &@              h@       @      V@      ,@                      @      1@              @      "@              7@      @      6@      @       @      @     �[@     @n@      @      3@      b@      ;@     �z@     @R@     `s@      b@      "@      @     �S@     @a@      �?      *@     @Y@      4@     �c@     �P@     �a@      Y@      @      @     �P@     �X@              $@      R@      ,@     �X@      J@     �Y@      R@      @              (@     �C@      �?      @      =@      @      M@      ,@     �D@      <@                      @@      Z@      @      @     �E@      @     �p@      @     �d@      F@       @              6@     �R@              @      :@      �?      i@      @     �^@      =@       @              $@      =@      @      �?      1@      @      Q@      �?      F@      .@              (@     `g@     �n@      (@      9@     Pq@     �J@     �r@     ``@     �s@      h@      4@       @      F@     �P@              @     @Q@      @     �Z@      4@     �W@     �J@               @      2@      *@               @      6@      @      @@      @      *@      (@               @      2@      &@               @      1@      �?      ,@       @      @       @                               @                      @       @      2@      �?      @      @                      :@     �J@              @     �G@      �?     �R@      1@     �T@     �D@                       @      A@              �?      8@      �?     �G@       @      ?@      8@                      2@      3@               @      7@              <@      "@     �I@      1@              $@     �a@     �f@      (@      4@      j@     �H@      h@     �[@     �k@     `a@      4@      @     �S@     �`@       @      (@      a@      <@      d@     �Q@     �c@      N@      *@      @     �Q@     �Y@      @      (@      _@      3@      a@     �K@     �`@     �H@       @               @      @@      @              (@      "@      8@      .@      8@      &@      @      @      P@     �G@      @       @      R@      5@      @@     �D@      P@     �S@      @      @     �@@      ?@      �?       @      L@      1@      1@      7@     �F@     �I@      �?       @      ?@      0@      @      @      0@      @      .@      2@      3@      <@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��<MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�8S��@�	           ��@       	                   �5@dI�"�@E           ��@                           �?g���G,@�           ̐@                           �?��#�غ@�            �@������������������������       �����I@�            �k@������������������������       ��l�}:'@9           �@                           �?A�	��@�            0u@������������������������       ��qH>s@C            �Z@������������������������       �+V�1S@�             m@
                           �?s���e	@�           ��@                          �:@��Wk�	@           ��@������������������������       ��5^��	@H           �~@������������������������       ��X~�o�	@�            �t@                           �?�5'ڍ�@�            �n@������������������������       ���k�~>@             �N@������������������������       ��ȳ�@r             g@                           �?S��@@           ��@                            �?�hgw�@g           ��@                           �?Wk�u���?R             `@������������������������       ���W�M�?.             R@������������������������       ���wfz9@$            �L@                           �?(���@           �{@������������������������       �3 �� @�            `p@������������������������       �;x����@r             g@                           @�*#��_@�           ��@                          �<@�0���@�           �@������������������������       ���7�{@�           Ѕ@������������������������       �F�z\��@            �C@                           @�:�q�@           �|@������������������������       �D��F@            �J@������������������������       ����0@�            Py@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     P�@      @@     �I@     `~@     �P@     ,�@     �h@     `�@     0v@      7@      .@      m@     �r@      7@      C@      v@      I@     w@     �d@     `v@     �k@      3@      �?     @V@     @`@      @      4@     @g@      .@     `o@     @R@      j@     �V@      @      �?     �S@      T@      @      2@     �`@      (@      b@      F@      b@     �Q@      @              >@      6@       @      @      7@      �?     �Q@      $@      I@      &@              �?      H@      M@      @      .@     @[@      &@     �R@      A@     �W@      N@      @              &@      I@      �?       @      K@      @     �Z@      =@      P@      3@                       @      $@                      .@              B@      @      @@       @                      @      D@      �?       @     �C@      @     �Q@      :@      @@      1@              ,@     �a@     �d@      1@      2@     �d@     �A@     �]@     �W@     �b@     �`@      ,@      ,@     �Z@     �`@      1@      1@     �`@      5@     @R@     �R@     �Z@     �[@      *@      @     �Q@      V@      (@      $@     �S@      &@      H@      G@     �R@      E@      @      &@     �B@      G@      @      @      L@      $@      9@      =@      ?@      Q@      @              B@     �@@              �?      ?@      ,@     �F@      3@     �E@      7@      �?              @      @                      @       @      7@      @      1@              �?              >@      =@              �?      ;@      (@      6@      .@      :@      7@                      U@      l@      "@      *@     �`@      1@     Є@      @@     `|@     �`@      @              8@     �U@      �?      @      >@      @      q@      &@      ^@      7@                              3@      �?              @      @     @R@      �?      1@       @                              @                      �?       @      I@              @      @                              (@      �?              @      �?      7@      �?      &@       @                      8@      Q@              @      7@      �?     �h@      $@     �Y@      .@                      &@      B@              @       @      �?     �`@      @      K@      $@                      *@      @@                      .@              P@      @     �H@      @                      N@     @a@       @      $@      Z@      *@     �x@      5@     �t@     @[@      @              >@     �U@      @      @      S@      $@     �n@      $@      j@     �L@                      <@      U@       @      @      N@      $@      n@      "@     �i@     �I@                       @      @       @      �?      0@              @      �?       @      @                      >@     �I@      @      @      <@      @     `b@      &@     @_@      J@      @              @       @               @      @              .@              @      1@      @              ;@     �H@      @      �?      8@      @     �`@      &@     �]@     �A@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�X�whG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @*Q���\@�	           ��@       	                   �3@�WdS��@|           T�@                           �?�����@�           `�@                           @v���@)           �}@������������������������       �MG?��@�            `x@������������������������       ��D��@7            �U@                            @�v��:@�            �m@������������������������       �S��&v�@j            �e@������������������������       �B�2l5�@*            @P@
                           �?��;��]	@�           x�@                           �?Q� �N�@           z@������������������������       �F�7{j	@�            �t@������������������������       �1��\�,@>            �U@                           �?B�5#�	@�           ��@������������������������       �H�H5�_@�            q@������������������������       ������	@�           `�@                           @�O� @+           |�@                           @����@�           ,�@                          �2@�����@�           ��@������������������������       ���
>1�?�            �z@������������������������       ��^��\�@�           x�@������������������������       �Ϝ��@             3@                          �5@2~fE�@M           ��@                          �3@�dp��|@�            Ps@������������������������       ���� q@t            @h@������������������������       �hﯳ@D            �\@                           �?'�0P��@�            �k@������������������������       ��N���@H            �\@������������������������       ��R�b@M            @[@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        5@     0q@     8�@      ?@     �Q@     `|@      R@     ȏ@     `m@     ��@     0w@      ?@      3@      i@     �s@      5@     �M@     �t@     �E@     �w@     �g@     Pw@      p@      ;@      @      G@     �W@      @       @     �V@      "@      g@     �I@     �b@     �Q@      @      @      ?@      O@      @      @     �Q@      "@      Z@      C@     @V@      L@      @       @      6@      I@      @      @      N@      @     �U@      6@      U@      H@              @      "@      (@                      $@       @      1@      0@      @       @      @              .@      @@              @      4@              T@      *@     �N@      .@                      *@      6@                      1@             �L@      @      H@      $@                       @      $@              @      @              7@      @      *@      @              *@     `c@      l@      2@     �I@     �m@      A@     �h@     `a@     �k@      g@      7@      �?     �D@     @P@      @      &@      O@      �?      T@      9@     �R@     �G@      @      �?      B@     �L@      @      "@     �I@              E@      5@      N@      F@      @              @       @               @      &@      �?      C@      @      ,@      @      �?      (@     �\@      d@      *@      D@      f@     �@@     @]@     �\@     �b@     @a@      2@              &@     �D@      @      &@      K@      @     �A@      2@      F@      F@      @      (@     �Y@     �]@      $@      =@     �^@      <@     �T@      X@     @Z@     �W@      &@       @     �R@      i@      $@      &@     @_@      =@     ��@     �F@     �{@     �\@      @       @      H@     @a@      �?      @     �S@      .@     0~@      9@     �r@     �P@      @       @      F@     @a@              @     @R@      *@      ~@      7@     �r@     @P@      @              @     �H@                      ,@             @k@      @     @Z@      9@               @     �B@     @V@              @     �M@      *@     �p@      0@      h@      D@      @              @              �?              @       @      �?       @       @      �?                      :@      O@      "@       @      G@      ,@      c@      4@      b@     �H@      �?               @      >@      @      @      6@      @      ^@      @     �U@      9@      �?              @      0@       @       @      0@             @S@      @     �N@      *@                      @      ,@      �?       @      @      @     �E@       @      9@      (@      �?              2@      @@      @      @      8@      $@     �@@      ,@      M@      8@                      $@      6@       @      @      ,@      @      2@      @      7@      (@                       @      $@      @      �?      $@      @      .@       @     �A@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@shzhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?3���iO@�	           ��@       	                    �?�*zu�5	@           ��@                           �?�tr�K@�           ��@                           �?R?�ԙ@}            �i@������������������������       �^�n��@9            @V@������������������������       �xC�{"@D            @]@                           �?��F��@           `|@������������������������       �H����@m            @f@������������������������       �<D�~@�            @q@
                          �7@ٿ���	@q           Ȏ@                           @i��rK�@^           h�@������������������������       �	B~#@�            �t@������������������������       �K�@�             l@                            @�C��0#
@           �z@������������������������       ��-0e�	@�            �m@������������������������       �YV�H�	@            �g@                            @������@�           ��@                          �4@k�eN/@�           ��@                            �?��ޗ j@p           �@������������������������       �St���@�           ��@������������������������       �ǳ��@�            pr@                          �7@��\�@!           �@������������������������       �I(�y��@            z@������������������������       �+ѬBT�@           �{@                           �?�Qr�@           �y@                          �1@�?��ҧ�?V            @^@������������������������       ���7~`u�?             >@������������������������       �0��f���?A            �V@                          �1@Uj�:@�            Pr@������������������������       ��W�_�0�?             B@������������������������       �7��!��@�            p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     P�@      5@      G@     @~@     @U@     ��@     �n@     ؇@     pu@      B@      (@      f@     �n@      .@      >@      p@      M@      l@     `c@     �o@     �g@      <@      @     �J@      Z@      @      $@     @\@      &@     �Z@     �O@     @\@     @Q@      "@      �?      :@     �B@                      ;@              C@      @      I@      5@       @      �?      @      (@                      2@              4@      @      8@      @                      5@      9@                      "@              2@      �?      :@      .@       @       @      ;@     �P@      @      $@     �U@      &@     @Q@     �M@     �O@      H@      @       @      "@      =@      @      @     �J@      @      9@      .@      3@      (@      @              2@      C@       @      @     �@@      @      F@      F@      F@      B@      @      "@     �^@     �a@      $@      4@      b@     �G@     �]@      W@     �a@     @^@      3@      @     �R@      S@       @      "@     �T@      ,@     @T@     �E@     �W@      P@      (@              H@     �D@       @       @     �B@      @     �O@      4@     �P@      B@      @      @      :@     �A@              �?      G@       @      2@      7@      =@      <@      @      @     �H@     @P@       @      &@      O@     �@@     �B@     �H@     �F@     �L@      @              A@     �A@      @      @      :@      4@      1@      :@      8@     �D@      @      @      .@      >@      @      @      B@      *@      4@      7@      5@      0@      �?       @     @^@     Pu@      @      0@     @l@      ;@     ��@      W@     �@      c@       @       @     �X@     @r@      @      ,@     �g@      9@     ��@      T@     `z@     �^@       @              B@     �d@       @      @     �R@       @      x@     �C@      k@     �O@      @              =@     �Y@       @       @      N@       @     pp@      7@     �c@      K@                      @      O@               @      .@             @^@      0@      N@      "@      @       @      O@      `@       @      $@     �\@      7@     �j@     �D@     �i@     �M@      @              C@     �O@      �?      @     �L@      $@      `@      &@     @T@      4@      @       @      8@     @P@      �?      @      M@      *@     @U@      >@      _@     �C@       @              7@     �H@       @       @      B@       @      e@      (@      V@      ?@                      �?      @              �?      @             �R@              =@      @                              @                                      6@              @                              �?      �?              �?      @             �J@              :@      @                      6@     �E@       @      �?      ?@       @     �W@      (@     �M@      ;@                      �?      @                                      3@              $@                              5@     �B@       @      �?      ?@       @     �R@      (@     �H@      ;@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��@p�*@�	           ��@       	                    �?��I׳�@�           z�@                            �?A�5�LR@�           ��@                           �?[hN��@�             x@������������������������       ������@�            p@������������������������       �W�x�ν@H            �_@                           �?ƺ��m@�            �s@������������������������       �k�j�@.            �R@������������������������       ���fy�@�            @n@
                           @{�FI}	@�           �@                           �?<s�d�
@�            �s@������������������������       ��a^� *
@�             m@������������������������       �2��3[@7            �T@                          �3@����.	@           �@������������������������       �c/�}@�            �w@������������������������       ��P�؆	@%           @�@                           �?�r	�o@8           0�@                          �3@E&���� @m           X�@                           @���$���?�            �r@������������������������       ��6�sn�?c            �e@������������������������       �DT���8 @X            @`@                          �5@���ߒ@�            �q@������������������������       �.��/w @H            @[@������������������������       �����@j             f@                          �1@N��T�@�           �@                           @1'���?�            `i@������������������������       ����̝��?U             a@������������������������       ��Y�䦄�?+            �P@                            @f�?Vmj@K           ��@������������������������       �=�욉@�           ��@������������������������       �t/'y��@f             d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     0q@     P�@      B@      K@     @{@      U@     <�@     �k@     ��@     �t@     �C@       @     �i@     `u@      ?@      E@     �r@      N@     px@      g@     px@     `n@     �B@             @Q@     �W@      @      @     �S@      @     `f@      =@     �d@      O@      "@              A@      H@      @       @      A@             �U@      *@     @]@      B@      "@              <@     �B@      @       @      :@             �G@      *@     �P@      ;@      @              @      &@                       @              D@              I@      "@      @             �A@      G@              @      F@      @      W@      0@     �H@      :@                      @      *@                      "@              ?@              *@       @                      =@     �@@              @     �A@      @     �N@      0@      B@      8@               @     @a@      o@      ;@     �A@     �k@     �L@     �j@     �c@      l@     �f@      <@      @      ?@     �I@      @      .@      I@      (@      5@     �@@     �H@     �A@      $@      @      =@     �A@      @      @      =@       @      *@      8@      D@      =@      $@               @      0@               @      5@      @       @      "@      "@      @              @     �Z@     �h@      5@      4@     �e@     �F@     �g@     �^@      f@     @b@      2@              9@     �L@      @       @      I@      $@     @Y@      ;@      N@      C@      @      @     �T@     �a@      0@      2@     �^@     �A@     �V@      X@      ]@      [@      (@       @      Q@     �j@      @      (@      a@      8@     @�@      B@     �{@     �V@       @              5@     �Q@              �?      ;@      @     `r@       @     �a@      1@      �?              &@      7@                      "@             �e@      @     �R@      "@      �?              @      *@                      �?             �Z@       @      D@      @                      @      $@                       @             @P@      �?      A@      @      �?              $@      H@              �?      2@      @     �^@      @     �P@       @                      @      4@              �?      @      �?     �K@      @      3@                              @      <@                      (@      @     �P@       @      H@       @               @     �G@     �a@      @      &@     @[@      2@      v@      <@     �r@     �R@      �?              �?      .@              �?      &@             @[@      @     �J@      "@                      �?      &@                      &@             �P@              E@      @                              @              �?                     �E@      @      &@      @               @      G@     �_@      @      $@     �X@      2@     �n@      8@     �n@     @P@      �?       @     �D@     @\@      @      @     @R@      1@     �i@      7@     �g@      J@                      @      *@      �?      @      9@      �?     �D@      �?      L@      *@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�B^dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�h';%P@�	           ��@       	                    @��W��@P           ֠@                           �?�u���@�           ��@                           �?dyT�b@�            �u@������������������������       �ҫ�iH @q            @f@������������������������       �]�Qst�@t            �e@                          �3@s����0@�            �@������������������������       �L�툃�@           0|@������������������������       �]���	�@�            p@
                           �?�.T��@�           $�@                           �?ӒH$���?            {@������������������������       ���X�?�             o@������������������������       ��nʊt�?p             g@                          �1@�JZP @�           ��@������������������������       ��P[`�x @w            �g@������������������������       ��m@0           �}@                           �?Y,/v��@Y           x�@                          �<@��o��@B           `@                          �;@2�q$�@            �x@������������������������       ����f�@@�            0w@������������������������       ��;^@             ;@                           @�pk(L@B             Z@������������������������       �����@1            @T@������������������������       ���K�� @             7@                          �?@1c��1	@           ��@                           @-}�E	@�           ��@������������������������       ���}f�	@�           �@������������������������       �]�.F�@           @z@                           @���4��@%            �P@������������������������       �x�^���@             ?@������������������������       �wR���@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     r@     ��@      B@     @P@     @@     �S@     8�@      g@     @�@     Pt@      ?@       @     @[@     pr@      3@      ?@     �l@      =@     ��@     �T@     0~@     �`@       @       @     �Q@     @c@      ,@      3@     �b@      6@     Pp@     �Q@     �i@     �T@      @              9@     �F@      @      @      @@      "@     �]@       @     �S@      9@                      (@      6@      @      @      2@      "@      O@      @      A@      @                      *@      7@                      ,@              L@      @     �F@      2@               @      G@     @[@      &@      *@      ]@      *@     �a@      O@     �_@      M@      @      @      <@      N@      @      @     �P@      @     �\@      D@     @S@      D@       @      @      2@     �H@      @      @     �H@      @      =@      6@     �H@      2@      �?              C@     �a@      @      (@     �T@      @      }@      (@     `q@      J@      @              &@      K@              @      .@             �n@      @     �U@      *@      �?              @     �@@              @      $@             �a@      �?     �E@      "@                      @      5@                      @             @Y@      @     �E@      @      �?              ;@     �U@      @      "@      Q@      @     �k@      @      h@     �C@      @              @      8@              @      &@             @R@      �?     �Q@      @                      8@     �O@      @      @     �L@      @     `b@      @     �^@     �@@      @      .@     �f@     pq@      1@      A@     �p@     �H@      q@     �Y@     Pt@     �g@      7@      @      G@     @T@              @      L@       @     �\@      1@      ^@      G@      @      @      A@     �N@              @     �F@       @      Z@      @      Z@      :@      @              >@     �J@              @      E@      @      Y@      @     @Y@      :@      @      @      @       @                      @       @      @              @                              (@      4@              @      &@              &@      $@      0@      4@      �?              (@      2@              @      $@                      "@      &@      1@      �?                       @                      �?              &@      �?      @      @              (@     �`@     �h@      1@      <@     �j@     �D@     �c@     �U@     �i@      b@      3@      @      ^@     @g@      0@      <@     �i@      D@     �c@     @T@     �h@     �`@      1@      @     �U@     �_@      &@      2@     �`@     �A@     �P@     @Q@     @Y@     �X@      1@              A@      N@      @      $@     @R@      @     �V@      (@      X@     �A@              @      ,@      (@      �?              @      �?       @      @       @      $@       @      @              @                      @      �?       @      @       @       @              �?      ,@      @      �?               @                       @      @       @       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{��GhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �7@��@x-�@�	           ��@       	                    �?(��t@�           ��@                           �?Kڝ��e@L           x�@                            �?��Èƨ@4           �~@������������������������       �K�ۮ(� @M            �`@������������������������       �3�j@�            `v@                            �?��-��@           @|@������������������������       ��? @T             `@������������������������       ����.@�            @t@
                          �1@C%LWE�@�           ��@                           @g�H倖@�            �w@������������������������       �2����@�            �u@������������������������       �ˣS���@             @@                           @9I�&u@�           Ė@������������������������       �)�r2/	@           ��@������������������������       ��<�((d@�           ��@                            �?�Ō��-	@�           ��@                           �?\'���@f           P�@                           �?���C�	@�            �q@������������������������       �$䍒�@K            �[@������������������������       �pJH@��	@m             f@                           @7O�h7@�            �p@������������������������       �CQo��=@w            �f@������������������������       �x%p~��@7            �U@                           @��;	@q           �@                          �?@�9��	@�            `x@������������������������       �BK�Q�	@�            0u@������������������������       �o��c�@            �I@                           @v�4�@z            �g@������������������������       ���U��J@l            @e@������������������������       �����|'@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     ��@      ;@      P@     @{@     �V@     p�@     @m@     X�@     �w@      A@      "@     �g@     0y@      (@     �F@     `r@      H@     (�@     @^@     8�@     �j@      6@              N@     �\@       @      @     �O@      @     px@      ;@     @k@     �H@      @              @@      P@              @     �C@      @     �j@      &@     @W@      7@      @              @      2@                      .@      �?     �P@       @      9@      @                      =@      G@              @      8@      @     @b@      "@      Q@      4@      @              <@     �I@       @              8@             `f@      0@     @_@      :@      �?               @      9@       @              @              F@      @      A@      @                      4@      :@                      2@             �`@      *@     �V@      4@      �?      "@     ``@      r@      $@      C@     �l@     �D@     �y@     �W@     �x@     �d@      2@              "@      I@      @      @      =@       @     �]@      5@     �Z@     �A@                      @      I@      @      @      8@              \@      1@     �Y@      =@                       @                       @      @       @      @      @      @      @              "@     �^@     �m@      @     �@@     @i@     �C@     pr@     @R@     0r@     ``@      2@      "@     �Q@      a@      @      :@     �`@      7@      \@      P@      ^@     @U@      (@             �I@     @Y@              @     @Q@      0@     �f@      "@     `e@      G@      @      $@     @[@     �a@      .@      3@     �a@     �E@      e@     @\@     �h@     �d@      (@      @     �H@     �P@      @       @     �N@      7@     �R@     �Q@     �X@     @V@       @      @      9@      @@      @      @      ?@      2@     �@@     �E@      A@     �J@      @       @      @      0@      �?              *@       @      8@      &@      0@      2@      �?      �?      2@      0@       @      @      2@      0@      "@      @@      2@     �A@      @              8@     �A@               @      >@      @      E@      ;@      P@      B@       @              1@      =@              �?      7@      @      <@      3@     �E@      .@       @              @      @              �?      @      �?      ,@       @      5@      5@              @      N@     @R@      (@      &@     @T@      4@     �W@     �E@     �X@      S@      @      @      J@     �J@      @       @     �M@      3@     �E@     �@@     �I@      K@      @      @      G@      J@      @      @     �H@      3@      E@      <@      F@     �C@      @      �?      @      �?       @      @      $@              �?      @      @      .@                       @      4@      @      @      6@      �?     �I@      $@     �G@      6@                      @      .@      @      @      1@      �?     �H@       @     �G@      6@                      @      @      �?              @               @       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ	��0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�Mc�n@�	           ��@       	                    �?m	Y��d@           x�@                           �?�ձ�@1            @                           �?L��M\@�             m@������������������������       ��;��@9             V@������������������������       ������@S             b@                          �8@�2��v@�            �p@������������������������       ���5�@{            �i@������������������������       �Bj��^@*             O@
                          �4@�*�`K@�           `�@                          �3@�
����?%           �|@������������������������       ��,|>v��?�            �w@������������������������       ��;z4��?8            �T@                           @�`]wX�@�            r@������������������������       �oZX{k�@�            @i@������������������������       ��y�@4            �U@                          �5@m�ђTl@�           ֤@                            @(��*�@�           �@                          �4@���Z��@�           x�@������������������������       ��-��@           ��@������������������������       ���f0\@x             h@                           �?���ٽ�@�            �v@������������������������       ��n�7S@             :@������������������������       �R��~�!@�            �t@                          �8@��<"�	@           ��@                           �?��(�@^            �@������������������������       �!dSj�l@�            �h@������������������������       �'.+@��@�            �u@                           @�֏��	@�            �@������������������������       ��g^�M2
@(           0}@������������������������       �X����A@�             n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     0t@     0�@      C@     �J@     pz@      W@     l�@     �l@     x�@     @x@      >@             �W@     �d@       @      &@     �U@      $@     �}@      F@     0p@     �X@      @             �P@      S@       @      $@      G@       @     @Y@      @@     @Z@     �K@      @              .@     �A@       @      @      7@       @      L@      1@      H@      ;@      �?              @      (@                      @             �B@      @      7@      @                      (@      7@       @      @      2@       @      3@      ,@      9@      6@      �?             �I@     �D@              @      7@             �F@      .@     �L@      <@       @             �@@      ;@               @      0@             �D@      (@     �I@      6@                      2@      ,@               @      @              @      @      @      @       @              =@     �V@              �?      D@       @     0w@      (@     @c@     �E@                      5@      C@              �?      5@             �p@      �?     �V@      7@                      3@      ?@                      (@             `j@             �T@      5@                       @      @              �?      "@             �J@      �?       @       @                       @      J@                      3@       @     �Z@      &@      P@      4@                       @      ?@                      "@      @     @U@       @     �F@      &@                              5@                      $@      @      6@      @      3@      "@              .@     �l@      v@      B@      E@     u@     �T@     �@     `g@     �~@      r@      ;@      @      U@     �j@      $@      5@     �b@      >@     0x@      Q@      s@     �`@      $@              O@     �d@      @      &@      [@      4@     �r@     �H@     @n@      W@      @             �L@      ^@      @      @     �U@      $@     �p@     �E@     �g@     �R@      @              @      F@              @      5@      $@      >@      @      J@      1@              @      6@     �I@      @      $@      D@      $@     @V@      3@      O@      E@      @              �?      @              @      �?      @       @      @       @       @              @      5@      F@      @      @     �C@      @     �U@      .@      N@      D@      @      &@      b@      a@      :@      5@     �g@      J@      h@     �]@     �g@     �c@      1@      @     @Q@      O@      &@      @     �W@      5@      [@      @@      S@     �J@      @       @      :@      <@      @       @     �A@       @     �E@      $@      6@      3@      @      �?     �E@      A@       @      @      N@      3@     @P@      6@      K@      A@               @     �R@     �R@      .@      ,@     �W@      ?@      U@     �U@      \@     �Y@      $@       @      F@      K@      &@       @     �J@      >@      F@     �R@      N@     �Q@      $@              ?@      5@      @      @     �D@      �?      D@      *@      J@      @@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJQ�XLhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?]S��ؠ@�	           ��@       	                    �?����	@�           ��@                           �?�Q���z@*           p}@                            @�5���@t            @f@������������������������       ������Q@Y            �a@������������������������       � ܓ;�� @             C@                          �5@(*��'F@�            Pr@������������������������       ��{�e�@Z             c@������������������������       ����PK+@\            �a@
                           �?��7��	@�           ��@                            @��'� �@           �y@������������������������       �LQx	�@�            0q@������������������������       �I�[�ߝ	@Z            �`@                           @|I�".
@�           x�@������������������������       ��W�3	�	@�           X�@������������������������       �h{]�+j	@>             Y@                           �?��;h�X@�           �@                            �?�WvM�@�           ��@                           �?C����9 @s            `h@������������������������       ��Uڷ���?;            �W@������������������������       �a`��@8            @Y@                           �?�4�<T�@U           ��@������������������������       ���z���@�            �s@������������������������       �.ضf@�            `n@                           @����R@�           T�@                           @'��|?#@           `|@������������������������       ��1��@�            �w@������������������������       �Э23<@,            �Q@                          �1@ ��V�@�           <�@������������������������       �� ��dW @}            �h@������������������������       ��CT@Y@F           @�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �t@     ؁@      C@     �I@      ~@     @V@     8�@      n@     X�@      v@      =@      1@     �g@     �l@      9@      @@     �n@     �N@      j@     �a@     �l@     `i@      5@              I@     �S@      �?      "@      M@      @     �W@      =@     �V@     �H@      @              3@      9@                      7@              C@      @      J@      0@       @              .@      2@                      5@              :@      @     �C@      0@       @              @      @                       @              (@              *@                              ?@      K@      �?      "@     �A@      @      L@      :@     �C@     �@@      @              0@      4@      �?       @      (@      @      G@      *@      2@      0@      @              .@      A@              @      7@      �?      $@      *@      5@      1@              1@     @a@     �b@      8@      7@     `g@      L@     �\@     �[@     @a@     @c@      .@       @      A@     �P@      @      &@     �R@      @     �L@     �A@      N@      J@      @      �?      1@     �F@      �?      @     �L@      @     �B@      >@     �D@      B@      �?      �?      1@      6@      @      @      2@      @      4@      @      3@      0@      @      .@      Z@     �T@      4@      (@      \@     �H@      M@      S@     �S@     �Y@      $@      "@     �X@     �Q@      3@      (@     �X@      F@     �C@     �M@      R@     �V@      @      @      @      *@      �?              *@      @      3@      1@      @      &@      @      �?     �a@     `u@      *@      3@     `m@      <@     ��@     @Y@     0�@     �b@       @              D@     @Z@      �?      �?      G@      @     @t@      8@     �f@      :@      @              �?      5@      �?              (@       @     �X@             �G@      "@      @                      @                      "@      �?      J@              6@      @                      �?      .@      �?              @      �?     �G@              9@      @      @             �C@      U@              �?      A@       @      l@      8@     �`@      1@      �?              1@     �F@              �?      :@       @     �b@      "@     @P@      @                      6@     �C@                       @             @S@      .@     �Q@      &@      �?      �?     �Y@     �m@      (@      2@     �g@      8@      y@     @S@      w@     �^@      @             �B@      W@      @      @     @S@      "@      T@      C@     @S@      B@                      9@     @R@      @      @      Q@      @     �R@      :@     �Q@      @@                      (@      3@                      "@      @      @      (@      @      @              �?     @P@      b@      "@      *@      \@      .@      t@     �C@     0r@     �U@      @               @      7@               @      @              W@      @     �L@      *@              �?     �O@     �^@      "@      &@     @Z@      .@     �l@      B@     @m@     �R@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ2�KDhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �1@�f+1v@�	           ��@       	                    @���N�@�            �@                           �?.ln�a@�            �r@                           �?���h @�            �m@������������������������       �X�>"@/            �R@������������������������       ��s���?u            `d@                           @�zK͒>@%            �O@������������������������       ���=��V@             >@������������������������       �|���#6�?            �@@
                           @�ֵ���@�            @s@                            @��g��@�             q@������������������������       �}� ��@�            �i@������������������������       ����=�@0             Q@                           @*��v�@             A@������������������������       �
1TUG@
             7@������������������������       ��t��`��?             &@                          �;@�P�x" @           ҩ@                           �?�?��@           P�@                           �?�=����@           (�@������������������������       ���h�j@�            �v@������������������������       �2L�re@<           �}@                           @[���lQ@�           ��@������������������������       ��5+K�@O           L�@������������������������       �:�!O��@�             q@                           @�hۑB�	@           |@                          �<@�� �	@�            �s@������������������������       ��Dd,(�	@/            �R@������������������������       ���*Ct	@�             n@                           �?%nm��B@O            �`@������������������������       ���|\�8@            �H@������������������������       �}���@3            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     `u@     `�@      @@     �I@      ~@     �V@     (�@     �k@     0�@     Pv@      8@              2@     �R@       @      @      D@      @     �p@      3@     �`@     �F@      �?              $@      ;@              �?      0@             `c@      *@     �N@      0@      �?              @      8@              �?      ,@             �^@      @     �K@      $@      �?               @      (@                      $@              <@      @      ,@      @                      @      (@              �?      @             �W@      �?     �D@      @      �?              @      @                       @             �@@      "@      @      @                      @      �?                       @              @      "@      @      @                               @                                      :@               @      @                       @      H@       @      @      8@      @      \@      @     @R@      =@                      @      G@       @       @      4@             �X@      @     �Q@      9@                       @     �A@              �?      0@              R@      �?     �N@      2@                      @      &@       @      �?      @              ;@      @      "@      @                       @       @              �?      @      @      *@       @      @      @                       @       @                      @      @      @       @      @       @                                              �?                       @                       @              3@     @t@     ~@      >@     �G@     �{@     �U@     І@     �i@      �@     �s@      7@      &@     �p@      z@      9@     �B@     `w@      O@     ��@      e@     X�@     `m@      3@              O@      Z@      �?      @      U@       @     `q@      @@     �i@     �K@      @              F@      M@      �?      @      H@       @     @Q@      2@     �V@      :@      @              2@      G@              �?      B@      @      j@      ,@      ]@      =@              &@     `i@     �s@      8@     �@@      r@      K@     �y@      a@     �u@     �f@      0@      @     �e@     Pp@      5@     �@@     p@      G@     �v@     @Y@     0t@     �b@      &@      @      ?@     �I@      @             �@@       @      G@      B@      :@      =@      @       @     �M@     @P@      @      $@     �P@      9@      E@     �A@     �J@     @S@      @       @      F@     �E@      @      $@      E@      8@      1@      >@      =@      N@      @      @      (@      .@      �?       @      $@      @      @      �?      @      "@      �?      @      @@      <@      @       @      @@      2@      &@      =@      7@     �I@      @              .@      6@      �?              8@      �?      9@      @      8@      1@                      @      $@                      @              0@      @      "@      @                      &@      (@      �?              5@      �?      "@       @      .@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ悠hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���G@�	           ��@       	                   �1@���\�@`           �@                           �?�+{I�@~           Ȃ@                           �?5�X���@s            �e@������������������������       ��ﾚ�@2            �Q@������������������������       �&�<?a@A            �Y@                          �0@M�g�+@           �z@������������������������       �~�0aL��?]            @b@������������������������       �W�_@�@�            �q@
                            @
���p@�           l�@                           @X��<4@�           �@������������������������       ��č�]6@E           `@������������������������       ��o��@�            �@                           �?�J�f�@            z@������������������������       �廤No@�             p@������������������������       �96�J2S@f            �c@                           �?�7�NE�@=           T�@                          �<@�|��@,           �}@                           �?�?�#
@�            Px@������������������������       �٠ֳ@u            @f@������������������������       �^`��@{            `j@                            �?;9����@<            @V@������������������������       �pdL�S�@             9@������������������������       ��.F��@,             P@                           �?01��J	@           ܓ@                            @��T��=
@@            �Y@������������������������       �o�\�	@&            @P@������������������������       �VՕ�M^@            �B@                           �?Rn;��@�           D�@������������������������       ���fGJ<
@c           ��@������������������������       �ZȠ�Ә@n           �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     0�@      =@      J@     |@     @T@     x�@     @k@     8�@     `v@      <@      @     �_@     �s@      @      5@      k@      A@     ��@     �X@     �~@     `e@      "@      �?      5@     @T@       @      @     �I@      �?     �k@      3@     @d@     �B@       @      �?      .@      8@       @       @      >@      �?      A@       @     �C@      0@                      @      &@                      1@              7@      @      &@      �?              �?      (@      *@       @       @      *@      �?      &@      @      <@      .@                      @     �L@               @      5@             @g@      &@     �^@      5@       @                      <@                      @              Q@      �?     �C@      @                      @      =@               @      2@             �]@      $@      U@      ,@       @      @     �Z@     @m@      @      1@     �d@     �@@      |@      T@     pt@     �`@      @      �?     �U@     �f@      @      *@      X@      5@     �t@      P@     �m@     �Y@      @      �?      J@     �N@       @      $@      O@      *@      W@      H@     �W@     �O@      @             �A@     �^@      �?      @      A@       @     `n@      0@     �a@     �C@      �?      @      3@     �I@       @      @     @Q@      (@     �\@      0@     �V@      @@      @      @      1@      8@      �?      @     �M@      $@      L@      $@      H@      8@       @               @      ;@      �?      �?      $@       @     �M@      @      E@       @      �?      *@     �g@     `m@      6@      ?@      m@     �G@     u@     �]@     �s@     `g@      3@      �?      F@     �P@      @      @     �M@      @      a@      ,@     �Y@     �C@      �?      �?     �A@     �K@      @       @      H@      @     @^@       @     �W@      .@      �?      �?      :@      @@      @       @      =@      �?      =@      @     �D@      @      �?              "@      7@                      3@      @      W@       @     �J@       @                      "@      &@              @      &@      �?      .@      @      "@      8@                      @      @                      @      �?      �?              @      @                      @      @              @      @              ,@      @      @      4@              (@      b@      e@      3@      :@     �e@      D@      i@     @Z@     �j@     �b@      2@      @      .@      @              @      .@      @      @      $@      1@      &@      "@      @       @      �?              @      @      @      @      @      ,@       @      @              @      @                       @      �?      �?      @      @      @      @      "@      `@     �d@      3@      3@     �c@      B@     `h@     �W@     �h@      a@      "@      "@     �M@     �W@      0@      .@     @R@      ;@     �L@      O@     �P@      R@      "@             �Q@     @Q@      @      @     �U@      "@     @a@     �@@     �`@     @P@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{k�+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?(j�IVa@�	           ��@       	                     �?�ߚ�ݐ@           P�@                          �>@I;5�@�           ��@                           �?�8,�`@�           �@������������������������       �WSA��]@�            Pu@������������������������       �t/�Ӆ@�            �r@                          �?@�Ъ��@             5@������������������������       ��	�o�� @             $@������������������������       �@	B0f@             &@
                           �?�TJ���@j           ��@                          �5@zT�(�|@�            Ps@������������������������       �!)?��}@v            �h@������������������������       �[~@G�P@K            @\@                          �3@��yP�@�            pp@������������������������       �-����@M             ]@������������������������       ��'��@\            `b@                          �4@��O@�           �@                           @�S!n��@�           8�@                           �?���@j           ��@������������������������       �f�WJ	@�            �w@������������������������       ��/�n@y            @g@                           @?'�x��@e           ��@������������������������       ������@W            `c@������������������������       �V����@           �{@                           @�t>���@�           ��@                           @HSh���	@\           �@������������������������       �͟�Cm�	@�            �j@������������������������       ��m�Yu	@�           h�@                           @�#{H6@o            �@������������������������       �@A���@`           �@������������������������       �*2�7�@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        =@      u@      �@      B@     �I@     �@     �S@     �@     `j@     `�@     �s@      =@             @X@     �c@      �?      $@     �_@      @     �{@      G@     q@     �Q@      @             �N@     @T@      �?      @     �Q@      �?      j@      6@     �d@     �D@      @              N@      S@      �?      @     �Q@              j@      ,@     �d@      C@      @              :@      C@      �?      @      E@             �`@      &@      N@      5@      @              A@      C@                      <@             @R@      @     �Z@      1@      @              �?      @              �?      �?      �?      �?       @              @                               @                      �?              �?      @               @                      �?      @              �?              �?              @              �?                      B@      S@              @      L@      @      m@      8@     �Z@      =@      �?              3@      F@              @      7@      @      a@      (@     �J@      *@                      &@      *@              �?      (@      @     @[@      "@      ;@      "@                       @      ?@              @      &@              ;@      @      :@      @                      1@      @@              �?     �@@             @X@      (@      K@      0@      �?              @      "@              �?      &@              M@      @      8@      @      �?              ,@      7@                      6@             �C@      "@      >@      $@              =@     �m@     pv@     �A@     �D@     �w@      R@     8�@     �d@     �@     �n@      6@      *@     @Q@     �c@      ,@      .@     �`@      .@      u@     �O@     �n@     �V@       @      *@     �C@     @T@      $@      "@      W@      &@     �]@      H@      V@      I@       @      *@      @@      D@      @      @      Q@      &@     @R@      ?@      O@      A@       @              @     �D@      @       @      8@              G@      1@      :@      0@                      >@     �S@      @      @      E@      @     `k@      .@     �c@     �D@                      ,@      9@                      (@      @      L@      @      8@      ,@                      0@     �J@      @      @      >@             `d@      "@     �`@      ;@              0@     @e@      i@      5@      :@     �n@     �L@     �n@     �Y@     @p@      c@      ,@      0@     �`@     @`@      .@      6@     �c@      I@     �V@     �T@     �_@      X@      $@       @      @@      7@      @       @      C@      1@      &@      4@      D@      (@      @       @     �Y@     �Z@      "@      4@     �]@     �@@     �S@     �O@     �U@      U@      @             �A@     �Q@      @      @     �V@      @     `c@      3@     �`@     �L@      @              =@     @Q@      @      @     @T@      @     �b@      ,@     �`@     �L@      @              @      �?       @              "@      @      @      @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����{Z@�	           ��@       	                    �?tc�*;*	@�           �@                           �?�Wi��@.           �}@                            @�X��@s             g@������������������������       ��j��,@S             `@������������������������       ���C9C @             �K@                           �?�����@�            r@������������������������       �
~P��@\            �a@������������������������       ���w���@_            `b@
                           �?�7T��	@�           ��@                           @B���@           �{@������������������������       �K|�hx@�            w@������������������������       �Y.JY�-@$            �R@                          �5@R�)�J
@�           h�@������������������������       �3ʍA��@�            q@������������������������       ��s[
@           �y@                          �7@0��q�N@�           �@                            @i�#x@0           ��@                            �?J����D@y           <�@������������������������       �:�2ڝ!@c           ��@������������������������       ��m�`L@           �{@                           @:5:���@�            0q@������������������������       �C���j�@�            �o@������������������������       ����鯆 @             7@                          �8@h�#a�@j           (�@                           �?�۹U��@S            �`@������������������������       �!�ρ=�@.             R@������������������������       �L0�T�@%             O@                            @ޔ�{@           �}@������������������������       �轗�}{@�            �v@������������������������       �Z�}���@D            @\@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     0s@     @�@      @@     �G@     @}@      U@     ��@      k@     ��@     �w@      @@      1@     `d@     �k@      7@      9@      p@     �E@     0p@     @a@      n@     �g@      :@              I@      O@       @      @      L@      @      `@      A@     �V@      D@       @              ,@      4@                      6@             �P@      @      E@      ,@                      &@      (@                      5@              C@      @      ?@      *@                      @       @                      �?              <@      @      &@      �?                      B@      E@       @      @      A@      @      O@      <@      H@      :@       @              $@      5@       @      @      *@      @     �B@      0@      8@      &@      �?              :@      5@               @      5@              9@      (@      8@      .@      �?      1@     @\@     �c@      5@      3@     @i@      D@     ``@      Z@     �b@     �b@      8@      �?      <@     �P@      @      &@     @U@      @     @T@      <@     @Q@      L@      @      �?      ,@     �K@      @      "@     @Q@      @      S@      9@      O@     �G@       @              ,@      (@               @      0@       @      @      @      @      "@      @      0@     @U@     �V@      1@       @     @]@     �@@      I@      S@     @T@     �W@      1@      @      ;@      C@               @     �K@      $@      9@      6@      G@     �A@      @      $@      M@     �J@      1@      @      O@      7@      9@      K@     �A@     �M@      $@      �?      b@     �t@      "@      6@     @j@     �D@     ��@     �S@     `�@     @g@      @             �V@     �p@       @      1@     ``@      ;@     ��@      D@     0v@     �_@      @             �T@     �k@      @      ,@     �\@      5@     ��@     �@@     �q@     �Z@       @              K@     �b@      @       @     �R@      1@     �v@      1@     �i@     @T@                      <@     �R@              @     �C@      @      f@      0@     �R@      9@       @               @     �F@      @      @      1@      @      V@      @     @R@      5@       @              @     �B@      @      @      .@      @     �U@      @      P@      5@                      �?       @                       @              �?              "@               @      �?      K@      P@      �?      @     �S@      ,@     �_@     �C@      e@     �M@       @      �?      *@      (@                      ;@      �?      @@      @      >@      &@       @      �?      @      @                      *@              0@       @      4@      @       @              @      @                      ,@      �?      0@      @      $@      @                     �D@      J@      �?      @      J@      *@     �W@      A@     `a@      H@                      A@      E@              @      F@      *@      M@      ;@     @\@      ?@                      @      $@      �?      �?       @              B@      @      :@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ1��ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�b�%}@�	           ��@       	                    �?��L�	@�           0�@                           �?���0�@,           @@                          �1@e�'��C@r            �g@������������������������       �	"���?            �C@������������������������       �XQc�3@Y            �b@                            �?Z7��g@�            �s@������������������������       �����l�@9             W@������������������������       ��UV�@�            �k@
                           �?��q19
@�           `�@                          �9@�@W�9o	@
           �y@������������������������       �]�NSh�@�            �s@������������������������       ���rŪ@:             W@                           @�	)�`
@�           �@������������������������       �C�:D�-
@�           ؂@������������������������       ���!�Ar	@?            �X@                           @w5	@�           ��@                           @�%�i@z           @�@                          �<@|ge�@j           P�@������������������������       ��ك�6�@D           `�@������������������������       ��8�̯@&             O@                            �?o!YO��@             >@������������������������       � �)7-@	             3@������������������������       ���^~@             &@                          �5@J�d �@/           T�@                           @B�R�2 @�           H�@������������������������       ����L@R           ��@������������������������       ��<(=�@�            �p@                           @����l@2           �~@������������������������       �?��@�            �o@������������������������       �jI#=@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     0s@      �@      8@     �Q@     �z@     @W@     h�@     �j@     X�@     v@      C@      6@      g@     `n@      *@     �G@     �j@     �J@      l@     �a@      p@     �g@      ;@      �?     �I@     �T@              "@     �P@      @     �[@      7@     �X@     �J@       @      �?      (@      9@                      5@              N@      @      H@      .@      �?                      �?                      @              7@              "@                      �?      (@      8@                      .@             �B@      @     �C@      .@      �?             �C@      M@              "@     �F@      @     �I@      2@      I@      C@      �?              $@      :@               @      @       @      0@      @      2@      "@                      =@      @@              @     �C@      �?     �A@      .@      @@      =@      �?      5@     �`@      d@      *@      C@     `b@      I@     @\@     @]@     �c@      a@      9@      @     �@@     �O@      @      4@     �K@      (@     �K@      D@      M@     �O@      @       @      <@     �K@      @      4@     �F@      @      H@      :@      G@      D@      �?      �?      @       @      �?              $@      @      @      ,@      (@      7@      @      2@      Y@     @X@      "@      2@      W@      C@      M@     @S@      Y@     �R@      4@      (@     @W@     @S@       @      2@     �S@     �A@     �G@     �N@     �W@     �P@      *@      @      @      4@      �?              ,@      @      &@      0@      @      @      @             �^@     s@      &@      8@     �j@      D@     h�@     �R@     X�@     `d@      &@             @Q@     �a@      @       @     @[@      @@     pq@      H@     �k@     �U@      @             �P@     �a@      �?       @     @Z@      9@     `q@      G@     �j@      U@      @             �L@     �`@      �?       @     �W@      9@     0q@      F@     �h@     �Q@       @              $@      @                      &@              @       @      ,@      *@       @               @              @              @      @      �?       @       @      @                                      @                      @      �?      �?      @      �?                       @                              @                      �?       @       @                      K@     �d@      @      0@      Z@       @     `@      ;@     �t@      S@      @              9@      [@       @      $@      H@      �?      w@      ,@     �g@      A@      @              1@     �R@       @      @      <@              q@      ,@      \@      ,@      @               @      A@              @      4@      �?     �X@             �S@      4@      @              =@     �L@      @      @      L@      @     �`@      *@      b@      E@      �?              2@      @@               @      <@             �T@      @     �P@      2@      �?              &@      9@      @      @      <@      @     �H@       @     �S@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��:EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@e�'��;@�	           ��@       	                    �?�"$BQ@�           �@                            @@�g�QE@�           X�@                           �?�/B4��@>           �~@������������������������       �.���� @�            Pp@������������������������       ����b�T@�            `l@                           �?��},��@c            `d@������������������������       �¬J!X�@2             T@������������������������       �>㷃1h@1            �T@
                           @]���@�           ܒ@                          �3@�x<�|j@�            �@������������������������       �ok\��@!           �}@������������������������       �d����@k            �d@                           @ȸ=���@o           ��@������������������������       ��D��=@R            �_@������������������������       �^��F�@           �{@                           �?�� Ar@*           �@                           �?��a �	@�           ��@                          �;@.�U&)
@�            �v@������������������������       ��;���	@�            @p@������������������������       ��f�3	@B            �Y@                           �?f)�	@�           0�@������������������������       ��s� 
�@^             b@������������������������       ��d>r	@7           `@                          �<@a���up@�           \�@                            �?||e_�"@W           ��@������������������������       �m_�%ѱ@�            �l@������������������������       ����Ok@�           ��@                            �?ga͚�@M            �^@������������������������       �:x9f�<@&             L@������������������������       �_���p@'            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      8@     @P@     �}@     �S@      �@     �j@     h�@     @u@      =@      @     @[@     �l@      "@      7@     �g@      6@     H�@      S@      y@     �a@      @              :@     �P@              @      G@      @     pr@      .@      c@     �C@      �?              2@     �J@              @     �A@             @l@      (@     �[@      =@      �?               @      7@              @      5@             �`@       @     �K@      ,@      �?              0@      >@                      ,@              W@      @      L@      .@                       @      ,@              �?      &@      @     @Q@      @      E@      $@                      @      @                      @      @      B@      �?      2@      @                      @      @              �?       @             �@@       @      8@      @              @     �T@      d@      "@      3@     �a@      1@      v@     �N@     �n@      Z@      @      @     �M@     �R@      "@      *@     �[@      (@     �`@      K@     �X@     �P@      @      @      I@      K@       @      @     @Q@      "@     �\@      F@     @Q@      J@       @       @      "@      5@      @      @     �D@      @      5@      $@      =@      ,@       @              8@     �U@              @     �@@      @     `k@      @     �b@      C@                      @      =@                      @      @     �E@      @      7@      $@                      1@     �L@              @      <@      �?      f@      �?     �_@      <@              .@     �g@     0s@      .@      E@     �q@     �L@     pw@     @a@     �y@     �h@      8@      (@     �]@      e@      .@      ?@     �b@      >@      ]@     �W@     �b@      [@      0@      @      D@      Q@       @      (@      H@      2@      D@     �D@      A@     �D@      @      �?      A@      H@      @      "@      A@      $@     �B@      7@      9@      ;@      @      @      @      4@       @      @      ,@       @      @      2@      "@      ,@              @     �S@      Y@      @      3@     @Y@      (@      S@     �J@     @]@     �P@      $@              1@      <@              �?      4@              6@      @      D@       @      @      @     �N@      R@      @      2@     @T@      (@      K@      I@     @S@     �M@      @      @     �Q@     `a@              &@     �`@      ;@     0p@      F@     `p@     @V@       @      @      N@     �^@              "@     @Z@      9@     �n@     �B@      n@     �Q@      @              0@      2@               @      =@      @     @T@      @     �L@      .@       @      @      F@     @Z@              @      S@      2@     �d@     �@@     �f@     �K@      @              $@      0@               @      >@       @      ,@      @      6@      3@      �?              @      @               @      &@      �?      @      @      ,@      $@      �?              @      &@                      3@      �?      &@       @       @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�7�EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@Q?���.@�	           ��@       	                     �?&���@p           �@                           @��۸�
@h           H�@                           �?�cv���@�            �r@������������������������       ���
@��@E            �Z@������������������������       ��+�<�@�             h@                           �?����}�?�            �o@������������������������       ��H���h @Q             `@������������������������       �0�Kغ��?Q            �_@
                           @��V"��@           ��@                           �?[��a�D@�           ��@������������������������       �&�ܦ��@�            �r@������������������������       �!xeS%�@1           �~@                           @���Td�@           H�@������������������������       �}�}�@x           ��@������������������������       ��'��t@�            �m@                           �?�F
4�@[            �@                           �?���ή

@$           ؊@                           �?�w=�!�@�             m@������������������������       � M����@-            �S@������������������������       ���)_@f            @c@                           @����y
@�           ��@������������������������       �$e��Qu
@�            �@������������������������       ��"��~@	             3@                          �7@���\?@7           (�@                          �6@*H��
�@�            pt@������������������������       ��*Y�}@q             g@������������������������       �{ϐ*��@`            �a@                           �?�B�ѝ�@f           ��@������������������������       ��v� 2�@\            @a@������������������������       ��Y�Gd�@
           @y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �q@     ��@      ?@     �I@     �z@     �X@     T�@      i@     8�@     �s@      A@      @      \@     �s@      (@      >@      h@      C@     ��@     �V@     `@      c@       @              4@     @U@               @      H@      "@     @h@      8@     `a@      >@       @              .@     �K@              �?     �B@      "@     �O@      7@     �S@      ,@       @               @      ;@                       @              5@      @      D@      @                      *@      <@              �?      =@      "@      E@      4@     �C@      "@       @              @      >@              �?      &@             ``@      �?      N@      0@                              ,@              �?      "@              K@             �B@      *@                      @      0@                       @             @S@      �?      7@      @              @      W@      m@      (@      <@      b@      =@     ��@     �P@     �v@     �^@      @      @      P@      \@      "@      4@      V@      6@     �f@      M@      c@      R@      @      @      :@     �E@      @      &@      >@      $@     �R@      9@      D@      A@               @      C@     @Q@      @      "@      M@      (@      [@     �@@     @\@      C@      @              <@      ^@      @       @      L@      @     �u@      "@     @j@     �I@      �?              3@     �S@      �?       @      9@      @      q@      @     �c@     �A@      �?              "@     �D@       @      @      ?@      �?      S@       @     �J@      0@              1@     `e@     �n@      3@      5@     @m@     �N@     t@     @[@     u@     �d@      :@      .@     �Z@     �^@      *@      2@      a@     �C@     @X@     @Q@     @^@     �X@      8@      �?      B@     �B@      @      @      C@      @      A@      $@     �D@      7@      �?      �?      &@      (@                      .@              5@      �?      (@      @                      9@      9@      @      @      7@      @      *@      "@      =@      2@      �?      ,@     �Q@     �U@      $@      *@     �X@      B@     �O@     �M@      T@     �R@      7@      *@      Q@     �U@      $@      *@     �V@      B@     �O@     �J@     �S@     �R@      5@      �?       @                              @                      @      �?               @       @     @P@      _@      @      @     �X@      6@      l@      D@      k@     �P@       @              <@      J@      @      �?     �G@      @      Z@      @     @Q@      0@                      2@      5@      @      �?     �@@      �?     �N@      �?     �A@      $@                      $@      ?@                      ,@      @     �E@       @      A@      @               @     �B@      R@      @       @     �I@      2@      ^@     �B@     `b@     �I@       @              @      ,@                       @       @     �G@      @     �J@      @      �?       @      ?@      M@      @       @     �H@      0@     @R@      ?@     �W@      F@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@[jc�0@�	           ��@       	                   �1@�]-F>@�           �@                           �?�jasi�@�           �@                           @����>@�             s@������������������������       �muk��s@�            �l@������������������������       ��ʞ�@,            �R@                            @Z'��@�            u@������������������������       �_��C��@�            �n@������������������������       ��bS5F@6             W@
                           �?8
OAY@           �@                           �?P�/cy@           �z@������������������������       � ���@p            `e@������������������������       �|/w��t@�            @p@                           @�Ú�*:@�           ��@������������������������       �p���^G@�            �u@������������������������       ���={�@           �{@                           �?qWbG�b@            �@                          �<@%���>�@o           ؁@                           �?��|�:@;            @������������������������       �R��3�@�            @q@������������������������       ��	��]q@�            �k@                           �?������@4            �R@������������������������       ���
Dm@             C@������������������������       �(ePg�@            �B@                           @I�79��@�            �@                          �:@�OQ$�	@J           Ȍ@������������������������       �G*2}	@�           H�@������������������������       �n�m� 	@�             q@                            �?'�	�>@g           x�@������������������������       ��T��/@�            �q@������������������������       ���fc�@�            q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@      r@     ��@     �@@      L@     �|@     @S@     l�@     �j@     p�@     pt@      B@       @     �Y@     �l@      &@      .@     `e@      4@     ��@      T@     0z@     �`@      *@       @      <@     @R@              @      J@             �q@      2@     �b@      @@      @       @      .@      @@              @      7@              b@      @      N@      1@                      &@      8@                      5@             �Y@      @     �L@      $@               @      @       @              @       @              E@      @      @      @                      *@     �D@                      =@             �`@      &@     �V@      .@      @              $@     �@@                      *@             �Y@      @      Q@       @      @              @       @                      0@              @@      @      6@      @              @     �R@     �c@      &@      (@     �]@      4@     �w@      O@     �p@     �Y@      $@      @     �C@     �C@      @       @     �P@      (@      U@      A@      U@     �I@      $@      @      $@      :@              �?      6@      �?      C@      ,@      A@      1@      @      @      =@      *@      @      �?     �F@      &@      G@      4@      I@      A@      @             �A@     �]@       @      $@      J@       @     pr@      <@      g@     �I@                      6@     @P@      @      @      =@       @     �W@      0@     @R@      <@                      *@     �J@      @      @      7@              i@      (@      \@      7@              @     �g@     �u@      6@     �D@     �q@     �L@     �x@     �`@     �v@      h@      7@              J@     @V@      @      "@     �P@      &@     �e@      1@     @\@     �A@                      G@      S@      @      @     �K@      $@     �d@      &@     �Y@      5@                      ;@      A@      @      @      8@       @     �[@      @      G@      (@                      3@      E@      �?              ?@       @      L@      @      L@      "@                      @      *@              @      (@      �?      @      @      &@      ,@                               @              @      @      �?      @      @      @      "@                      @      @              �?      @              @      @      @      @              @      a@      p@      1@      @@     �k@      G@     `k@      ]@     @o@     �c@      7@      @     �X@     �f@      .@      8@     �`@     �B@      V@     @X@     @\@     @Z@      5@      @     @R@     `a@      &@      5@     �Y@      ;@      N@     �O@      U@     �G@      1@      @      :@     �E@      @      @      >@      $@      <@      A@      =@      M@      @             �B@     �R@       @       @     �U@      "@     ``@      3@      a@     �J@       @              7@     �G@              @      8@      @     �P@       @     �R@      >@      �?              ,@      ;@       @      @     �O@       @     @P@      &@      O@      7@      �?�t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�>�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�i���1@�	           ��@       	                    �?�1�}XI@}           8�@                          �3@�~j���@�           Ȅ@                            �?m5�\@b           ��@������������������������       ��@��5 @\             c@������������������������       �����@           `z@                           �?��� r@A            �V@������������������������       ���W�<n@             =@������������������������       ��%^��@+             O@
                           @p�~8n@�           ԑ@                          �0@��v�j@t           �@������������������������       ����|��@             M@������������������������       �k�S��@V           @�@                           @+��]�@f           ��@������������������������       ���[�!@�            �v@������������������������       �|Σ0Ӣ@y            �h@                            �?�l�?KQ@:           v�@                           @���NV�@�           D�@                           �?�!�x9@i           ��@������������������������       �6^N.Z�@�            `s@������������������������       ��{���@�           ؄@                           @"VdS{	@S             `@������������������������       �B��H��	@=             U@������������������������       ���U��+@             F@                           �?K:���@~           P�@                           @����@�            �r@������������������������       ��Ս��%@t            �g@������������������������       �X�X��@C             [@                          �6@����v@�           �@������������������������       �ް���@�            �k@������������������������       ��+�̦9	@:           @~@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     ��@      ;@     �N@     �{@     �T@     �@      k@     �@     �t@      <@      @      Y@      p@      @      8@      e@      4@     �@     �V@     �v@      `@      @              C@      V@              @      G@              r@      3@     `a@      C@                     �@@     �Q@               @     �C@             `o@      0@     �_@     �A@                      @      :@                       @             @Q@      @      D@      @                      <@     �F@               @     �B@             �f@      (@     �U@      =@                      @      1@              @      @             �C@      @      (@      @                      �?      @                      �?              "@      @      @       @                      @      $@              @      @              >@              @      �?              @      O@     @e@      @      1@     �^@      4@     �u@     �Q@      l@     �V@      @      @     �D@     �U@      @      &@     �S@      ,@     �[@     �O@     @Z@      K@      @               @      5@              �?      @              ,@              "@       @              @     �C@     �P@      @      $@      S@      ,@      X@     �O@      X@      G@      @              5@     �T@      �?      @      F@      @     �m@       @      ^@     �B@                      1@      J@              @      E@      @     �a@      @      U@      3@                      @      ?@      �?      @       @       @     �W@      @      B@      2@              $@     `i@     �s@      5@     �B@     0q@      O@     @x@     �_@     p{@     �i@      8@      @     �[@     �d@      @      ;@     �`@     �D@     �f@      T@     �l@     @[@      ,@      @      W@     �c@      @      :@      ^@     �@@      e@     �K@      j@     �Y@       @      �?      :@      J@       @      @     �C@      @     �Q@      @     �Q@      ?@      @      @     �P@      Z@      �?      6@     @T@      <@     �X@      I@      a@     �Q@      @      �?      2@      &@      @      �?      *@       @      (@      9@      7@      @      @      �?      (@      &@      @      �?      $@      @      @      2@       @      @      @              @                              @      @       @      @      .@       @              @     @W@     �b@      .@      $@     �a@      5@     �i@     �G@      j@     �W@      $@              =@     �I@      �?      �?      @@       @     �V@      *@      O@      .@                      8@      B@      �?      �?      7@       @      F@      &@      B@      $@                      @      .@                      "@              G@       @      :@      @              @      P@     �X@      ,@      "@     �[@      3@     @]@      A@     @b@      T@      $@      �?      2@      :@       @              D@      @     �B@      @      Q@      4@       @      @      G@     @R@      (@      "@     �Q@      0@      T@      =@     �S@      N@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{��<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @a���Q@	           ��@       	                    �?Kϕ�@N           �@                            �?T� �.@�           �@                           �?ig����@x            �i@������������������������       �y�8�3@S             `@������������������������       �r��`��@%            @S@                            �?��ܴD@           P{@������������������������       �_�Qs1@[            �b@������������������������       ��QUY*�@�             r@
                           �?o���p	@�           �@                          �2@��Lk��@           @z@������������������������       ���R��@8            �V@������������������������       ��Gha��@�            �t@                           !@�gwzջ	@�           ��@������������������������       ��F���	@�           @�@������������������������       �I �D�J@             1@                           �?�O���#@1           �@                          �3@e�����@n           H�@                            �?�|J1o�?�             s@������������������������       �z�m^���?*             P@������������������������       ����yw�?�             n@                          �8@�I[���@�            �q@������������������������       ��0��*@z            @i@������������������������       ���P�׿@3            �S@                           @e���:@�           �@                          �<@�+ێ�@�           ��@������������������������       �h����@�           ��@������������������������       �lPTJP�@"            @P@                          �6@�14�{�@             8@������������������������       ���!zȓ@             "@������������������������       ��3����?	             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �r@     (�@      ?@      H@     �z@     �U@     ��@     `j@     Љ@     0v@      ?@      6@     @k@     �u@      7@      ?@      r@     �P@     �v@     @f@     0x@     �l@      :@       @      P@     @X@      @      @      P@       @     �c@      =@     �d@     �H@      @       @      2@      D@              @      (@              F@      @     �P@      *@      @       @      *@     �A@              @      @              1@      @      C@      $@      �?              @      @                      @              ;@              <@      @      @              G@     �L@      @      @      J@       @      \@      :@     �X@      B@      �?              @      1@       @       @      *@              B@      *@     �C@      3@      �?             �C@      D@      �?       @     �C@       @      S@      *@     �M@      1@              4@     @c@     @o@      4@      8@     @l@     @P@     �i@     �b@     �k@     �f@      5@       @      ?@     �S@              (@     @Q@      @     �Q@      :@      N@     �N@      @       @      &@      ,@                      @              5@      &@      (@      (@                      4@      P@              (@      O@      @      I@      .@      H@     �H@      @      2@     �^@     �e@      4@      (@     �c@     �M@      a@     �^@     `d@     @^@      1@      2@     �^@      e@      4@      (@     `c@     �K@      a@     �^@     `d@      ^@      (@              �?      @                       @      @              �?              �?      @      @     �S@     @m@       @      1@     �a@      4@     ��@     �@@     p{@      _@      @              4@      S@      �?      @     �@@      @     0q@      "@     �`@      ;@      �?              "@      >@              �?      @              f@      @     @P@       @      �?                      �?                      @             �E@              ,@      @                      "@      =@              �?      @             �`@      @     �I@      @      �?              &@      G@      �?      @      :@      @     �X@      @     @Q@      3@                      &@      B@      �?      @      2@      �?     �S@      �?      F@      "@                              $@                       @      @      4@       @      9@      $@              @     �M@     �c@      @      *@     �Z@      .@     v@      8@     s@     @X@      @      @      J@     �c@      @      &@      Y@      .@     �u@      6@     �r@     @X@      @      @      F@     �a@      @      &@     �U@      .@     �u@      6@     `r@     @T@      @               @      .@      �?              ,@               @              "@      0@                      @      �?      �?       @      @               @       @       @                                              �?       @      @              �?               @                              @      �?                      @              �?       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�eLhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��a@�	           ��@       	                    �?L��j9�@v           �@                           �?�?7oR@�           ��@                          �3@�tL�,�@�             x@������������������������       ��5dg�K@�            0q@������������������������       ��(O^c@G            @[@                           @�ڴ��@�            @w@������������������������       �r%%K,@z             g@������������������������       ��2?ѐ�?p            `g@
                           @8�(	��@�            �@                           @�ʕr@�           Ї@������������������������       �����@G           �~@������������������������       ��8(|Z@�            �p@                           @C�6E��@�           0�@������������������������       �+�z��	@j             d@������������������������       ����\L�@>           `~@                           �?�����@9           T�@                          �:@3S�K�	@           ��@                          �7@��|2�@=           p�@������������������������       ��nʛ�P@�            @p@������������������������       ��,����@�            �p@                           @*�S��m
@�            �t@������������������������       ������"
@�            Pr@������������������������       �$B�-�@            �D@                          �7@"Ce��%@%           ȋ@                           �?$sa�P>@�            `s@������������������������       �	��#[@/            @S@������������������������       �_}�؋�@�             m@                           �?��F�@i           �@������������������������       ��u�s[@_            �a@������������������������       ��,��@
           p{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �r@     ��@      >@      M@     �~@      U@     8�@      i@     P�@     �v@      <@      @     �]@     Ps@      $@      :@     �l@      >@      �@     @T@      ~@      d@       @             �G@     �X@               @     �J@       @     `t@      .@      f@     �A@      �?              1@      J@              �?     �@@       @      e@      (@     �S@      4@                      (@      =@                      5@      �?     �]@      $@      Q@      0@                      @      7@              �?      (@      �?     �I@       @      $@      @                      >@     �G@              �?      4@             �c@      @     �X@      .@      �?              3@      9@              �?      0@             �I@      �?     �N@      &@                      &@      6@                      @             �Z@       @     �B@      @      �?      @     �Q@     @j@      $@      8@      f@      <@     �w@     �P@      s@     �_@      @      @      H@     @^@      "@      1@      ^@      3@     �b@     �L@     @^@      V@      @      @      ?@      O@      @      &@     �U@      0@     �V@      @@      W@     @P@              @      1@     �M@      @      @      A@      @     �M@      9@      =@      7@      @              7@     @V@      �?      @     �L@      "@     �l@      "@     �f@      C@       @               @      8@                      *@      "@      K@      @     �A@      (@       @              .@     @P@      �?      @      F@             �e@      @     �b@      :@              1@     �f@     �o@      4@      @@     @p@      K@     pr@     �]@     �r@     �h@      4@      .@     �X@     �a@      .@      7@     �b@      <@     @U@     �S@     �[@     �X@      2@      �?     �R@      V@      @      2@      Y@      &@     �I@     �H@     @R@      G@       @      �?     �G@      F@       @      &@      F@      @      ,@      2@      D@      @@      @              ;@      F@      @      @      L@      @     �B@      ?@     �@@      ,@      @      ,@      9@      K@       @      @      H@      1@      A@      =@     �B@     �J@      $@       @      7@     �I@       @      @      E@      .@      ?@      1@      B@      H@      "@      @       @      @                      @       @      @      (@      �?      @      �?       @     �T@     �[@      @      "@      \@      :@     @j@     �D@     �g@      Y@       @              E@     �C@       @      @     �F@      �?     �W@       @      H@     �@@                      @       @       @              "@              B@              $@       @                      C@      ?@              @      B@      �?      M@       @      C@      9@               @     �D@      R@      @      @     �P@      9@      ]@     �C@     �a@     �P@       @              @      3@                      @       @      I@      @      D@      @               @      C@     �J@      @      @      N@      1@     �P@      @@      Y@     �N@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�F+��@�	           ��@       	                    �?p�tX@�@�           t�@                          �6@� ���@�           ��@                           @� 5@           �|@������������������������       ���~���@�            p@������������������������       ���;G���?~             i@                           @Y��R*�@            �h@������������������������       �D�m�@`             c@������������������������       ��8�߱f @            �G@
                           �?�:��L@i           `�@                          �<@Ɲ��P@�             p@������������������������       �|���JW@�             l@������������������������       �B��9�g@             @@                            �?�� @�            �t@������������������������       ��\���3 @n            �f@������������������������       �̲hy���?a            �b@                           @�h����@�           ؤ@                          �4@i��^w�@�           |�@                           �?�b�y@�           x�@������������������������       �.ڢ���@-            @Q@������������������������       ���%c	@w           Ȏ@                            �?�����@E           ��@������������������������       �؋_o��@�            �v@������������������������       ��w;`@a           ��@                           !@վߘL	@�            �r@                          �7@bk�(8	@�            �q@������������������������       ��*fhw@i             c@������������������������       �� ~?�@V            �`@������������������������       �η:@
             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@      r@     �@      1@     �A@     �|@     �U@     P�@     @j@     ��@     u@      8@             �K@     �d@       @      @     �[@      (@     �{@     �F@     �t@     �Q@      �?              :@     �Q@       @      @     �Q@      (@     �p@      :@     �a@     �A@                      $@      I@              �?     �F@      $@     �j@      4@      X@      ,@                      $@      7@                      ?@      $@      Y@      0@     �L@      $@                              ;@              �?      ,@              \@      @     �C@      @                      0@      5@       @       @      9@       @     �M@      @     �F@      5@                      (@      0@       @       @      9@      �?      C@      @      @@      5@                      @      @                              �?      5@      @      *@                              =@      X@              @     �D@              f@      3@     �g@     �A@      �?              4@      L@              @      =@             �G@      (@     �P@      6@                      3@     �H@                      9@             �F@      $@      P@      (@                      �?      @              @      @               @       @      @      $@                      "@      D@                      (@              `@      @     @^@      *@      �?              @      >@                      @              K@       @     �S@      @                      @      $@                      @             �R@      @      E@       @      �?      2@     `m@     �y@      .@      =@      v@     �R@     X�@     �d@     X�@     �p@      7@      *@      i@     �v@      *@      <@     0s@      L@      �@     �`@     �}@     �n@      .@      @     @S@      e@      @      @      Z@      @     `t@     �H@     �l@     �S@       @       @      @      "@              �?      *@       @      @      @      0@       @               @     �Q@     �c@      @      @     �V@      @     �s@      F@     �j@     �Q@       @      "@      _@     `h@       @      7@     `i@     �H@     �g@      U@     �n@     �d@      *@      @      E@      P@              $@     �J@      3@      F@      <@      N@      B@      @      @     �T@     ``@       @      *@     �b@      >@     @b@      L@     `g@     ``@      $@      @      A@      H@       @      �?     �F@      3@     �C@      @@      H@      5@       @      @      @@      F@       @      �?     �E@      *@     �C@      @@     �G@      5@      @              &@      ;@      �?      �?      <@      @      <@      ,@      4@      ,@      @      @      5@      1@      �?              .@       @      &@      2@      ;@      @       @               @      @                       @      @                      �?              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��%�M@�	           ��@       	                   �;@�1OW	@�           �@                           �?��*y	@^           �@                           �?�N�%@           �x@������������������������       ��MW?1.@{            �h@������������������������       �I9ڗC�@�            `h@                           �?%d��{�	@]           ��@������������������������       ��x�6�	@�            �s@������������������������       ���FO�	@�           ��@
                           @�UW}	@�            �o@                          �?@���Ԫ'	@�             l@������������������������       �����D@m             e@������������������������       �e֍�Q?@!            �L@                          �=@���	\�@             >@������������������������       �EA��W�?             *@������������������������       ���1�@             1@                           @33���@�           �@                           @v��|�@�           ��@                          �3@���4S|@�           ��@������������������������       ���{�O/@�            �m@������������������������       ��2�C@�            Pv@                          �7@lJ�w�@�            �x@������������������������       �����?@�            r@������������������������       ��J��&�@?             Z@                          �6@�O
���@8           ̔@                          �4@��3LZ�@O           �@������������������������       ����Z;@�           �@������������������������       �y��r@�             l@                           @�5&��@�             w@������������������������       �� ���?@�            �u@������������������������       ����(��@
             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ?@     r@     �@      9@      L@     �|@     @U@     ��@     �i@     ؈@     �u@      ;@      =@      e@      q@      5@     �@@     �l@      F@     `j@     @]@     �o@     �g@      7@      .@     �`@     @m@      4@      =@     �i@      @@      h@     �Y@     @k@     �a@      2@              <@     @R@       @      @      K@       @      U@      7@     @W@      <@       @              0@      ?@       @      @      =@       @      D@      0@     �E@      ,@      �?              (@      E@                      9@              F@      @      I@      ,@      �?      .@      Z@      d@      2@      :@      c@      >@      [@     �S@     @_@     @\@      0@      @      @@     �P@      &@      @      J@      $@      :@      3@      =@      I@      @      "@      R@     �W@      @      3@      Y@      4@     �T@      N@      X@     �O@      "@      ,@     �B@      D@      �?      @      8@      (@      3@      .@      A@      I@      @      (@      B@      A@      �?      @      6@      $@      &@      (@      A@     �F@      @      @      7@      9@              �?      0@      $@      $@      @      >@      C@      @      @      *@      "@      �?      @      @              �?      @      @      @               @      �?      @                       @       @       @      @              @      �?                                                       @      @       @              @               @      �?      @                       @               @      �?               @      �?       @      ^@     �r@      @      7@      m@     �D@     �@     �U@     ��@     �c@      @       @      P@     �c@              (@     @]@      ;@     �q@     �F@      j@     �R@      �?             �E@      U@               @     �S@      .@     `b@      C@     ``@     �I@                      &@      E@              @      2@              S@      (@      N@      .@                      @@      E@              @      N@      .@     �Q@      :@     �Q@      B@               @      5@      R@              @     �C@      (@     �`@      @     @S@      7@      �?              ,@      L@                      2@      (@     @\@      @     �M@      *@      �?       @      @      0@              @      5@              6@      @      2@      $@                      L@     `b@      @      &@     �\@      ,@     @�@      E@     �t@      U@      @              =@     �[@      @      @      T@      @     �z@      @      o@      G@      @              9@      S@      @      @     �H@             0v@      @     `f@      C@       @              @      A@              �?      ?@      @      R@             @Q@       @      �?              ;@     �B@      �?      @     �A@      $@     @W@     �A@     �U@      C@                      4@     �A@      �?      @     �@@      @      W@      ?@     �U@      C@                      @       @                       @      @      �?      @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJmehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�g��o @�	           ��@       	                   �7@�~���'@           $�@                           @���Cn@D           ��@                          �1@����,@           `z@������������������������       ��~V�@C            �[@������������������������       �2�wzU@�            �s@                          �5@xa�D @8           �@������������������������       �3�BO��?           �{@������������������������       �D	�Q�� @)            �O@
                            @^ҭ��@�            �r@                           �?w��ǄA@�             j@������������������������       ��@���@@             Y@������������������������       ��j��6�@C             [@                           �?Hk��9�@<            �V@������������������������       �+�R0@%             M@������������������������       ���B��@            �@@                           @��:��@�            �@                           �?u��,/	@�           ��@                           @k<���q	@�           T�@������������������������       �N��6f	@k           ��@������������������������       �~,���P@W            �_@                           �?�iR��@           �y@������������������������       �	��k	�@             @@������������������������       �M�>@�            �w@                          �7@����ݻ@�           H�@                          �4@�T�@�@           ��@������������������������       �r�z7?@a            �@������������������������       ���jK��@�            q@                           @�wA* `@�            �s@������������������������       ��3��T�@v            �f@������������������������       �}����@U            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      q@     h�@      ;@     �F@     `}@     �R@     ��@     �l@     ��@     �t@      :@             �S@     �e@       @       @     �Z@      "@     �|@     �B@     Pq@     �Q@      @             �J@     �]@       @       @     @Q@       @     �x@      3@     �j@     �H@                      C@      I@      �?             �C@      �?     �`@      3@      ]@      :@                      @      "@                      2@             �I@      @      1@      @                      ?@     �D@      �?              5@      �?     @T@      .@     �X@      6@                      .@     @Q@      �?       @      >@      �?     �p@             @X@      7@                      .@      K@               @      ;@      �?     �m@             @V@      ,@                              .@      �?              @              ;@               @      "@                      :@     �J@              @     �B@      @      N@      2@      P@      5@      @              ,@      G@              @      1@      @      A@      *@      J@      .@      @              "@      7@               @      @      @      5@      @      4@      &@                      @      7@              �?      *@      @      *@      @      @@      @      @              (@      @              @      4@              :@      @      (@      @                      @      @              @      *@              *@      @      &@      @                      @      @                      @              *@       @      �?      �?              3@     `h@     x@      9@     �B@     �v@     �P@     Ȃ@     �g@     H�@     �p@      3@      2@     �a@     �l@      *@      ?@     �o@      L@     @m@      c@     �h@      f@      0@      2@      Z@     �c@      *@      8@     �i@     �C@      b@     @[@     `a@     `a@      .@      0@      X@      b@      *@      8@      f@     �@@      a@     �S@     �`@     �^@      &@       @       @      *@                      >@      @      "@      ?@      @      1@      @              B@     �R@              @     �F@      1@     @V@      F@      M@      C@      �?              @      @              @      @                      @      @      @                     �@@     �P@               @     �D@      1@     @V@      D@     �K@      @@      �?      �?     �K@     @c@      (@      @      \@      $@     �v@      C@     @t@      V@      @              ;@     @^@      @      @     @P@      @     �s@      ,@      n@      K@       @              0@     �R@      @       @     �@@      @     @n@      ,@     �c@      B@                      &@      G@       @       @      @@      @      R@             @U@      2@       @      �?      <@     �@@      @       @     �G@      @     �J@      8@     �T@      A@      �?      �?      0@      2@               @     �A@             �C@      @     �G@      2@      �?              (@      .@      @              (@      @      ,@      2@      B@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��PRhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�<��2@�	           ��@       	                     �?�X�?^�@�           \�@                           �?�n+��@�           ��@                          �<@-`*�e)	@�           (�@������������������������       �Ծ����@�           x�@������������������������       �����w�@C            �]@                          �<@��R�@�            �u@������������������������       �^3�m�@�            �t@������������������������       �.Q���"@             2@
                           �?bѱ�>~@�           0�@                          �<@��;@�            `r@������������������������       �����@�            @p@������������������������       ����Rgs@             A@                          �3@��u�k�@�           0�@������������������������       ���G-{%@�            �l@������������������������       �v��R	@d           ��@                          �4@;�}�@6           l�@                           �?T�`�@;           (�@                           @��Bl��@(           @}@������������������������       �,��c4 @�            �u@������������������������       �����Ǎ@N             _@                          �1@pB�P� @           {@������������������������       ���`���?c            �b@������������������������       �WuL��@�            �q@                           �?�O�)@�           ��@                            �?���åN@�            `x@������������������������       ���5`F@�            �k@������������������������       �x�6��@l             e@                          �9@�A�9�y@            y@������������������������       �{+���@�             q@������������������������       ��'_ Q@X            �_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     @q@     P�@      :@      I@     �}@      X@     �@     �j@     �@     �u@      =@      (@     �i@     �t@      3@      A@     u@     �S@     �v@      f@     z@     @l@      8@       @     @[@     @d@      $@      7@     @c@      E@     �f@     �V@     `l@      Z@      .@       @      T@     @Z@      "@      .@      \@      >@     �\@     �S@     ``@      U@      *@       @      R@     �V@      "@      *@     @X@      7@      Y@     �M@      _@      K@      &@               @      ,@               @      .@      @      ,@      3@      @      >@       @              =@     �L@      �?       @      E@      (@     @Q@      *@      X@      4@       @              <@     �K@      �?      @     �D@      $@     @Q@      $@     �W@      0@      �?              �?       @               @      �?       @              @       @      @      �?      $@     @X@     �d@      "@      &@     �f@     �B@     `f@     �U@     �g@     �^@      "@              8@      A@      �?      @      E@       @     @R@      5@      Q@      9@                      7@      >@      �?      �?      <@       @     @Q@      3@     �P@      5@                      �?      @              @      ,@              @       @       @      @              $@     @R@     �`@       @      @     �a@     �A@     �Z@     @P@     �^@     @X@      "@      �?      @      A@      �?       @      G@      @      M@      *@     �D@      8@              "@     �P@     �X@      @      @     �W@      ?@      H@      J@     @T@     @R@      "@       @     �Q@      l@      @      0@     �a@      1@     Ȃ@      C@     |@     �]@      @              <@      \@       @      "@      I@       @     �y@      "@      m@     �G@      �?              0@     �H@       @      @      =@             �j@      @      \@      B@                      (@      @@                      3@             `e@      @     �U@      5@                      @      1@       @      @      $@              F@       @      :@      .@                      (@     �O@              @      5@       @     @h@      @      ^@      &@      �?               @      ,@                      @              S@       @      H@       @      �?              $@     �H@              @      1@       @     �]@       @      R@      "@               @      E@     @\@      @      @      W@      .@      h@      =@      k@      R@      @       @      6@      O@      �?      @      J@      "@     @Y@      @     �U@     �C@      @              .@      B@               @      ;@      "@     �O@      @      J@      .@               @      @      :@      �?      @      9@              C@      @     �A@      8@      @              4@     �I@      @       @      D@      @     �V@      6@     @`@     �@@      �?              $@      F@                      7@       @      R@      ,@     �W@      ,@      �?              $@      @      @       @      1@      @      3@       @      B@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�phG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���}B_@�	           ��@       	                    �?��\���@\           �@                           �?�w�;�F	@�           ��@                          �6@�)h�e)@*           @|@������������������������       �Ν7ξ@�            �q@������������������������       �%bD��i@u            `e@                           �?""�P�	@�           ��@������������������������       �D�i���@           �y@������������������������       ����l^�	@�           �@
                            �?0ru�`�@l           H�@                           �?�"���@�            �u@������������������������       �MY�Ս�@A            @[@������������������������       �Y(z�@�            @n@                            @nL�(��@�            �p@������������������������       �ӣHG-@8            �S@������������������������       ��:�Q��@d            `g@                          �4@u,]7�@I           �@                           �?�V�@R           ��@                           �?\�7�V�?�             w@������������������������       �1u[����?�            �i@������������������������       ��o��?l             d@                           @�!���@a           8�@������������������������       �*$b�	@T            �`@������������������������       ���7@            z@                          �7@���s3�@�            �@                           @fz.9�q@�             y@������������������������       �g��@;            �W@������������������������       �{���8}@�            s@                          �<@1�<�N,@�            @y@������������������������       ����}X�@�             s@������������������������       �dNu�@?             Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     �@      =@     �P@     Pz@     @U@     �@     `k@     ��@     �x@      ;@      1@     �m@      s@      8@     �H@     �r@     �O@     �v@     `f@     �v@     �p@      4@      1@     @f@     �j@      4@      A@     �k@     �G@     �l@     �`@     �o@      j@      3@              G@     �N@       @      @     �I@      @     @Y@      <@     �V@      M@      @              <@      B@      �?       @      7@      @      V@      3@      L@      9@                      2@      9@      �?      @      <@              *@      "@     �A@     �@@      @      1@     �`@     �b@      2@      <@     `e@      F@      `@     @Z@     @d@     �b@      ,@      @     �B@     �M@      @      ,@     �Q@      ,@      Q@      A@     �P@      F@      @      ,@     �W@      W@      .@      ,@     @Y@      >@      N@     �Q@      X@     �Z@      &@             �N@      W@      @      .@     �R@      0@     �`@      G@     @\@     �M@      �?             �C@     �K@      �?      (@      C@      .@     @R@      7@     �Q@      8@      �?              ,@      (@               @      @             �B@       @     �@@      @                      9@     �E@      �?      $@     �@@      .@      B@      5@     �B@      4@      �?              6@     �B@      @      @     �B@      �?      O@      7@     �E@     �A@                       @      @                      4@              1@      "@      ,@      @                      ,@      ?@      @      @      1@      �?     �F@      ,@      =@      >@              �?     �S@     �i@      @      2@      _@      6@     ؄@      D@     �z@     �_@      @             �C@     @Z@       @      (@      E@      @     0{@      *@     @j@      M@                      &@      <@              @      (@              k@      @      R@      3@                      @      *@              @      @              `@       @     �@@      (@                      @      .@                      @             �U@      @     �C@      @                      <@     @S@       @      @      >@      @     `k@       @     @a@     �C@                      "@     �@@                      @      @      E@      @      <@      $@                      3@      F@       @      @      9@              f@      @     �[@      =@              �?      D@     �X@      @      @     �T@      3@      m@      ;@     �k@      Q@      @              .@      L@       @      @     �@@      &@     �`@       @     �Y@      B@      @              @      "@      �?               @       @     �@@              3@       @      @              $@     �G@      �?      @      9@      @     �Y@       @      U@      <@              �?      9@     �E@      �?      @     �H@       @     @X@      9@     @]@      @@      @      �?      *@      A@              @      ;@      @      S@      7@     �X@      3@      @              (@      "@      �?              6@      �?      5@       @      3@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�^�AhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @4�W2@�	           ��@       	                    �?ڪ�0��@o           0�@                           �?���k@�           ��@                            @vrGa�@%           �|@������������������������       �I��G@�            `o@������������������������       �Cjh@�            �j@                           �?�_7n�=@o            @d@������������������������       �����Oo@=            @W@������������������������       ��ʊ��@2            @Q@
                          �:@��ӵ[	@�           ��@                          �4@��kG"�@#           �@������������������������       ��.��@o           ��@������������������������       ���UX	@�           ��@                           �?��>7
@�            �r@������������������������       �e'&>[@-            �R@������������������������       ��|���

@�             l@                           �?�2�&�@(           Ě@                            @��{� @\           ��@                          �4@ �΀�� @#           �}@������������������������       �]�v�4�?�            @q@������������������������       �Y]{��@x            `i@                           @z8QU
��?9             V@������������������������       �I�y��?             B@������������������������       ���M�?"             J@                           �?[�D[�@�           �@                          �4@g��w2d@W           H�@������������������������       �Bc��@�            @p@������������������������       ���@�@�            Pp@                           @��YV�F@u           ��@������������������������       �G%����@f           Ђ@������������������������       �LSks�z@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      r@      �@      6@      J@      ~@     �S@     �@      k@     ��@      u@      >@      7@      j@     �u@      2@     �D@     �t@     @P@     �w@      f@      v@      m@      7@       @     @P@     @V@      @      @      T@      @     �d@      ;@      `@      J@      @       @     �G@     �S@      @      @     �N@      @     �Y@      5@     �W@      F@      �?       @      :@      A@      �?              D@             �F@      (@      N@      >@      �?              5@     �F@       @      @      5@      @      M@      "@      A@      ,@                      2@      $@              �?      3@      �?      O@      @     �A@       @       @               @      @              �?      ,@              D@      @      ,@      @                      $@      @                      @      �?      6@      �?      5@      @       @      5@     �a@     �o@      .@     �A@     �o@     �N@     �j@     �b@      l@     �f@      4@      &@      [@     �k@      $@      :@     �j@      F@     �h@     @\@     @h@     �^@      0@      "@      @@      W@      @      "@      V@      "@     �\@      H@     @Y@      P@      @       @      S@      `@      @      1@      _@     �A@     @U@     @P@     @W@     �M@      (@      $@     �A@     �A@      @      "@      E@      1@      0@     �B@      ?@      M@      @      �?      @      @      �?      @      5@              @      $@      "@      .@      �?      "@      ?@      ?@      @      @      5@      1@      &@      ;@      6@     �E@      @      �?      T@     �m@      @      &@     @b@      ,@     �@     �C@     �z@     �Y@      @              .@     @P@               @      ?@      �?     �p@       @     �b@      9@      �?              ,@      O@                      9@      �?     �k@       @     @_@      7@      �?              @      <@                      (@              d@      @     �L@      (@      �?              &@      A@                      *@      �?      N@      @      Q@      &@                      �?      @               @      @             �H@              9@       @                              @                                      6@              &@                              �?                       @      @              ;@              ,@       @              �?     @P@     `e@      @      "@     �\@      *@     @w@      ?@     �q@     �S@      @      �?      @@     �R@      @      @      O@      @      c@      "@      `@     �E@      @              *@      <@       @      @      8@             �W@       @     �P@      4@              �?      3@     �G@      �?       @      C@      @      M@      �?      O@      7@      @             �@@      X@      �?      @     �J@      "@     `k@      6@      c@     �A@      �?              :@     �W@      �?      @     �H@       @      k@      3@     �b@     �A@      �?              @      �?                      @      �?      @      @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJūyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�YC�W@�	           ��@       	                    �?���1�/@           ��@                           �?��R�/�@$           �|@                           �?5��<@i            �c@������������������������       �-r���@5            �U@������������������������       �T<Ի[�@4            �Q@                            �?����ì@�            s@������������������������       ��Hy�˰@=            @Y@������������������������       ��`I6a@~            �i@
                           �?x��K��@�           ��@                          �8@�A/��@           P{@������������������������       ����BHC@�            �v@������������������������       ���4�@*            �R@                            �?��\d@�            v@������������������������       ���Wq�@@z            �h@������������������������       �U��&z�?\            @c@                           @6^>�@�           Ȥ@                           �?�YK*�@�           :�@                          �8@�B��	@t           ��@������������������������       ��
��`�@�           �@������������������������       ��7�/

@�            �s@                           @*�-(�H@T           �@������������������������       �{B���@�            Pq@������������������������       ���o��@�           ��@                          �5@����@�            pt@                           @,G��	@X            �b@������������������������       ��g�G�	@9            �X@������������������������       ���2}�a@             I@                           @_圝#�@j            `f@������������������������       �?_��y@T            �a@������������������������       �SvoTm8@             C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     ��@      B@      J@      {@     @Q@     `�@     @j@     �@     �u@      <@       @      U@     �e@      @       @     �Y@      @     0|@     �B@     �s@      Q@      @       @      I@      R@      @      @     �J@       @     �Y@      9@      Z@     �D@       @       @      *@      5@                      *@             �G@      @      G@      $@               @      @      @                      "@              >@      @      8@      @                      @      ,@                      @              1@      @      6@      @                     �B@     �I@      @      @      D@       @     �K@      3@      M@      ?@       @               @      7@              �?      $@              6@      @      ;@      @                      =@      <@      @      @      >@       @     �@@      *@      ?@      ;@       @              A@      Y@      �?      @     �H@      @     �u@      (@      j@      ;@      �?              2@      J@              @      A@      @      j@      @     �V@      7@                      1@      C@              @     �@@      @     `f@             @R@      0@                      �?      ,@                      �?              =@      @      2@      @                      0@      H@      �?              .@       @     �a@       @     @]@      @      �?              "@      C@      �?              @       @     �P@      @     �Q@      @      �?              @      $@                      &@             �R@      @      G@      �?              0@      i@     �x@      =@      F@     �t@      O@     H�@     �e@     (�@     �q@      9@      ,@      e@     �u@      =@      E@     �q@     �D@     �@     �b@     `@     �m@      .@      *@     �X@     @a@      8@      ;@      c@      9@     �Z@     �W@     �c@     @a@      (@      @     @P@     @W@      (@      8@     �]@      .@     @T@     �G@     �^@     �U@      @      "@     �@@     �F@      (@      @      A@      $@      9@      H@      B@      J@      @      �?     �Q@      j@      @      .@     �`@      0@     �x@      K@     pu@      Y@      @      �?      0@     �K@      �?       @      @@      @      N@      8@      L@      4@                      K@      c@      @      @      Y@      (@      u@      >@     �q@      T@      @       @     �@@      I@               @     �G@      5@     �H@      8@     �G@      E@      $@       @      $@      1@               @      1@      .@      <@      @      4@      9@      @       @       @      (@               @      .@      .@      $@      @      @      0@      @               @      @                       @              2@              *@      "@      �?              7@     �@@                      >@      @      5@      3@      ;@      1@      @              4@      <@                      .@      @      3@      (@      8@      1@       @              @      @                      .@       @       @      @      @              �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�+fzhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@���5@�	           ��@       	                    �?��/��@�           ��@                           @�q`�4 @O           h�@                            �?	�@!@�             o@������������������������       ��1ԤT�@0            �R@������������������������       ���`�@o            �e@                          �2@�� *��?�            @q@������������������������       �'�5�w��?�            �k@������������������������       ��;<N���?!            �J@
                          �1@*���]�@F           �@                           @����~@�            �v@������������������������       ��@T"��@a            �c@������������������������       ��0o��=�?�            �i@                           �?��l�]�@e           ȁ@������������������������       �~��X\�@            �G@������������������������       ��~�ߒ�@F           P�@                          �:@���t>@           4�@                           @��	gQ�@�           ��@                           @�w�,@z           �@������������������������       ��'e�@           8�@������������������������       ��W�B:@v           ؂@                           @_�%��@.           ~@������������������������       ��V���R@�            s@������������������������       ��[߶@t             f@                          �<@���]y�	@n           ��@                          �;@������@�             n@������������������������       � ^|D�@X             `@������������������������       ��>�^Z�@E             \@                          �A@Q����u	@�            pt@������������������������       ��,*	@�            �s@������������������������       ��tc��@             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      r@     @�@      C@      H@     �z@     @S@     ؎@      j@     ��@      v@      :@      @     �R@     `h@      @      @      a@      0@     �@     �M@     @u@      Z@      @              8@     �M@               @     �B@      @      m@      &@     �`@      6@      �?              1@      :@                      ;@      @      T@      $@     �Q@      0@                      �?      *@                      @              3@      @      ;@      @                      0@      *@                      6@      @     �N@      @     �E@      &@                      @     �@@               @      $@              c@      �?      P@      @      �?              @      >@               @      "@              `@      �?     �E@      @      �?              �?      @                      �?              8@              5@      @              @     �I@      a@      @      @      Y@      *@     @q@      H@     �i@     �T@      @      �?      3@     �N@       @       @      1@      �?      _@      .@     �V@      <@              �?      0@     �A@       @      �?      $@      �?      A@      *@      6@      5@                      @      :@              �?      @             �V@       @     @Q@      @              @      @@     �R@      @      �?     �T@      (@      c@     �@@     �\@      K@      @       @              *@                      @      �?       @      @      ,@      @               @      @@      O@      @      �?     �S@      &@     �b@      =@     @Y@      H@      @      2@     �j@     Px@      @@     �E@     `r@     �N@     �}@     �b@     �@     @o@      5@      @     �b@     �r@      6@      ?@     `k@     �E@     �y@     @Y@     �z@     @d@      1@      @     �[@     `j@      *@      4@     @d@     �@@     �t@      I@      u@      _@      0@      @     �U@     @_@      *@      0@      ]@      ;@      `@     �E@     �b@     @U@      ,@      �?      7@     �U@              @      G@      @     �h@      @     �g@     �C@       @             �D@      W@      "@      &@     �L@      $@     �T@     �I@     @V@      C@      �?              ;@     �P@      @      &@      @@      @     �A@     �F@      J@      8@      �?              ,@      :@      @              9@      @     �G@      @     �B@      ,@              *@      O@     �U@      $@      (@     �R@      2@     @Q@      H@     �T@      V@      @      "@      7@     �B@      @       @      @@      @     �E@      8@     �B@      8@                      (@      6@       @              2@      @      5@      4@      ,@      0@              "@      &@      .@       @       @      ,@       @      6@      @      7@       @              @     �C@     �H@      @      $@     �E@      *@      :@      8@     �F@      P@      @             �B@     �H@      @      $@     �D@      *@      :@      7@      F@     �O@      @      @       @                               @                      �?      �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ=�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @(�D�7B@�	           ��@       	                    �?s����@e           ��@                           �?��Scb�@�           ��@                          �<@���g@7           ~@������������������������       �M���@           p{@������������������������       �>4��h�@             E@                            �?�mӱ	@l             f@������������������������       �d.U�,@&             L@������������������������       ��z���v@F             ^@
                           @��pb	@�           ��@                           �?��f�(	@N           t�@������������������������       �8b�!3�@I            �[@������������������������       �Vu��@           ��@                           @�Ẽ��	@t            �i@������������������������       ���S�x�@U            �b@������������������������       �{M|��V@            �K@                          �4@x���!�@A           <�@                          �0@�W�x��@R           ��@                           @<Ok�Q��?R            �_@������������������������       ���B]w'�?,            �Q@������������������������       �fcYI��?&            �K@                           �?�D|�V@             �@������������������������       �����c�?�             r@������������������������       �O "�@F           ��@                           @�$8m�@�           ��@                          �=@'����@�           ��@������������������������       �x'��v@�           X�@������������������������       ��Jޱ�@            �H@                           �?������@6            @U@������������������������       ��v?�q�@            �@@������������������������       �o�G��@"             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     ��@      =@     �H@     �z@     @X@     �@     `l@     X�@     v@     �A@      *@     �j@      u@      6@      @@     �q@     @R@     Pv@     �g@      x@     �l@      >@             @R@     �W@       @      @     �O@      @      c@      F@     @d@     �F@       @              L@      T@       @      @      J@      @     @W@      B@      [@     �D@      @              I@     @R@       @      @      G@      @     @W@      >@     �Y@      @@      @              @      @               @      @                      @      @      "@                      1@      .@               @      &@       @      N@       @      K@      @      @               @      @               @      @              0@              6@              @              .@      "@                      @       @      F@       @      @@      @              *@     �a@     `n@      4@      9@     �k@      Q@     �i@     `b@      l@      g@      6@      $@     �_@     �i@      4@      2@     �h@      M@      g@     �[@     �i@      d@      ,@      @      *@      $@              @      7@       @      @      (@      2@      1@       @      @     @\@     `h@      4@      (@      f@      L@     �f@     �X@     `g@     �a@      (@      @      0@      C@              @      5@      $@      4@     �B@      3@      9@       @      �?      (@     �@@              @      &@       @      2@      9@      $@      6@       @       @      @      @                      $@       @       @      (@      "@      @      @      �?     @Q@     �k@      @      1@      b@      8@     �@      B@     �z@     �^@      @              C@     �Z@              "@      J@      @     �{@      3@     `l@     �M@      �?              @      ,@                                      Q@              @@      "@                      @      @                                     �E@              5@                                      $@                                      9@              &@      "@                     �A@     @W@              "@      J@      @     `w@      3@     `h@      I@      �?              $@      6@               @      *@             �e@      @      M@      @      �?              9@     �Q@              @     �C@      @      i@      ,@      a@     �F@              �?      ?@     �\@      @       @     @W@      4@     `l@      1@     �h@      P@      @      �?      8@      Y@      @       @     �S@      1@     �i@      "@     �g@      N@       @      �?      3@     �X@      @      @      P@      1@      i@       @     �f@      I@       @              @      �?       @      @      .@              @      �?      @      $@                      @      .@       @              ,@      @      4@       @      $@      @       @              �?      @                      @      @      $@      @       @               @              @      "@       @              "@              $@      @       @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�i#ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�bF`B@�	           ��@       	                    �?GJ�$ޖ@}           r�@                           �?r_R�u�@�           p�@                          �;@2����@4           p~@������������������������       ���W�@	           z@������������������������       ���&��@+            �Q@                          �9@���֤@q            �d@������������������������       ��ׇWk�@^             a@������������������������       ��qՠ� @             ?@
                           �?��g0	@�           ��@                          �4@���~�*	@�           $�@������������������������       �thP��_@	           �z@������������������������       �Eu�eܭ	@�           ��@                           �?y~��/@            z@������������������������       ����~SB@             C@������������������������       ����W�@�            �w@                           @��	]\S@-           @�@                           �?"�\�_�@            �@                          �3@���L�@\           ��@������������������������       �H���  @�            r@������������������������       �+4Tځ�@�            �n@                           �?%<��@�           H�@������������������������       ������@�            �u@������������������������       �-a�@�            �t@                          �7@��t�G@            }@                          �4@����@�            0u@������������������������       �\�?6@�            �m@������������������������       �*��2�k@:            �Y@                            �?�bA@Q            @_@������������������������       �r�v(@#             M@������������������������       ��C��'�@.            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     ��@      <@     �C@     �}@     �S@     �@     �l@     ��@     Pz@      5@      3@      k@     Ps@      7@      @@     �t@      N@     �w@     �e@     �w@     �r@      .@      @     @P@     �V@               @     �R@      @     �d@      <@     �a@     �P@      @      @      H@     �Q@              @      M@       @     �Z@      ;@     @Z@     �L@       @              C@     @P@              @     �H@       @     �Y@      7@     �W@      B@       @      @      $@      @              @      "@              @      @      $@      5@                      1@      4@              �?      1@      @     �L@      �?      C@      $@      �?              .@      .@              �?      $@      @      K@              ;@      "@                       @      @                      @              @      �?      &@      �?      �?      0@      c@     @k@      7@      8@     p@     �J@     �j@      b@     �m@     �l@      (@      0@      ]@      e@      3@      0@     �h@     �C@     �`@     @Y@      d@     �f@      &@      @      ?@     �I@      @      @     @T@      �?     �Q@     �B@     @Q@     �R@              (@     @U@     �]@      ,@      &@     �]@      C@      O@      P@     �V@      [@      &@              B@     �H@      @       @      M@      ,@     @T@     �E@      S@      H@      �?              "@       @              @      �?      �?       @      @       @       @                      ;@     �G@      @       @     �L@      *@     �S@      B@     �R@      D@      �?      @     �S@     �k@      @      @     �a@      2@      �@      L@     �{@     �^@      @      @     �G@     �e@              @     �X@      1@     @{@      @@     �t@     �Q@       @              0@     �S@              �?      @@      @     �l@      "@     �`@      >@       @              $@      A@                       @             `a@      @     @T@      &@       @              @     �F@              �?      8@      @     �V@      @      J@      3@              @      ?@     �W@              @     �P@      *@     �i@      7@     �h@      D@              @      3@     �J@              @     �C@      �?     �W@      "@     @Y@      5@                      (@     �D@                      <@      (@      \@      ,@      X@      3@                      @@      H@      @             �D@      �?      b@      8@      \@     �J@      @              3@      F@      @              5@      �?      _@       @     �T@      @@      @              $@      ;@      @              (@             @V@       @     �O@      7@                      "@      1@                      "@      �?     �A@              4@      "@      @              *@      @      �?              4@              4@      0@      =@      5@      �?              @      �?                      @              @      $@      7@      "@                      @      @      �?              0@              0@      @      @      (@      �?�t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�8`�/@�	           ��@       	                   �<@��%��@U           ��@                          �5@��9_�@�           ؝@                           �?.���@�           �@������������������������       ������@�             y@������������������������       ����^"@�           ��@                           �?���TX	@           ��@������������������������       ��27l�@�            �k@������������������������       ��
�	@}           ��@
                            @Ee�h+�@�            �l@                           �?R����f@W             `@������������������������       ���Ҕ@             C@������������������������       �	ccT�@>            �V@                          �?@U�~p�O@;             Y@������������������������       ���	|Z @+            �P@������������������������       �RG>@            �@@                           �?���@F           ��@                           @J�"�� @�           ��@                           @�q��R�?�             y@������������������������       �)��J�_ @X            �b@������������������������       � �A�=z�?�             o@                           �?��@�            �l@������������������������       �Լ�H�M@K            @_@������������������������       �ĝ+�2�@C             Z@                           @��jl@�           �@                          �1@�u�7@�           T�@������������������������       �x/���?�             k@������������������������       �)&��@/           �@                          �4@-T��9�@            �B@������������������������       ��P��i�?             *@������������������������       ��nǤ�@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     `s@     �@      ?@     �J@     �{@      W@     h�@      j@     �@     �u@      ?@      (@     `j@     ps@      5@     �C@     s@     @S@     @v@     �d@     0y@     �j@      9@      (@     �f@     �q@      3@      =@     @p@     �O@     �u@     �b@     �w@     @e@      5@      @     �Q@     `e@      &@      ,@     �b@      ;@     @l@     @R@      n@     �X@      @      @      0@      R@      @      @     �P@      ,@     �U@      @@     �O@     �A@      @      �?     �K@     �X@      @      $@     @T@      *@     `a@     �D@      f@      P@      @       @     @[@     @[@       @      .@      \@      B@     �^@     �R@     �a@     �Q@      ,@       @      B@      ?@               @      5@      @      I@      @      K@      (@      @      @     @R@     �S@       @      *@     �V@      ?@      R@     @Q@     �U@     �M@      $@              ?@      ?@       @      $@     �F@      ,@       @      2@      7@      E@      @              1@      *@                      6@      $@      @      &@      .@      @@      @              @      @                       @      @              @      @      "@                      &@      @                      4@      @      @      @      &@      7@      @              ,@      2@       @      $@      7@      @      @      @       @      $@                      &@      1@       @      @      $@      @      @      @       @       @                      @      �?              @      *@                       @      @       @                     �X@     `i@      $@      ,@     �a@      .@     H�@      E@      }@     �`@      @              1@      Q@      �?              <@      @     �s@      $@     �c@      ?@      �?              "@     �E@                      ,@       @     �l@      @     @U@      ,@                      @      5@                      @       @     �R@             �A@      @                      @      6@                       @             �c@      @      I@      @                       @      9@      �?              ,@       @     �T@      @     �Q@      1@      �?              @      1@                      @       @      J@       @      @@      @                       @       @      �?              @              ?@      @     �C@      $@      �?             �T@     �`@      "@      ,@      \@      &@      u@      @@     @s@     �Y@      @             @S@     �`@       @      ,@     @Y@       @     �t@      @@     �r@      X@      @               @      4@                      "@              X@      @     �Q@      .@                     �R@     @\@       @      ,@      W@       @     �m@      =@      m@     @T@      @              @       @      �?              &@      @      @              @      @                              �?                                      @              @      @                      @      �?      �?              &@      @      �?               @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�|��,@�	           ��@       	                     @؀vEN�@           <�@                           �?�0���@B           0�@                          �;@�+��lD@4           �}@������������������������       ��2�2y�@           p{@������������������������       ����b�@             D@                          �6@���3�|@           pz@������������������������       �f�G�@�            `p@������������������������       ��j�`O@a             d@
                           �?쬪s	@�            �t@                           �? 7�F@}            �f@������������������������       �,biz�@?            �U@������������������������       �v���o�@>            �W@                           �?�����?`            �b@������������������������       ���9r\@6            @U@������������������������       �&���2�?*            �O@                          �4@i�D�@�           ��@                           �?Ai���7@�           <�@                           @����Œ@3            �U@������������������������       ��n�bQ@             L@������������������������       �Ꭿ���@             ?@                           @2��)�@�           ��@������������������������       ���H�ʝ@�            �@������������������������       ��ҍ�w�@           �y@                          �9@��7��@�           ��@                            �?�x�c@U           �@������������������������       ���.V�w@�             r@������������������������       �8��&�@�           �@                           �?9�VqlX	@V           P�@������������������������       �CY���	@�            �t@������������������������       �w{Gh�g@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     @s@     ��@      ?@     �F@     �|@     @S@     ��@     `l@     ��@     �u@      :@      �?      T@     �e@      @      &@     @^@      1@     �{@     �C@     q@     �O@      @      �?      N@     �`@       @      @     @T@      1@     �s@      9@     @k@      H@      @      �?      =@     �P@      �?       @      G@      $@     �g@      (@      W@      =@      �?              ;@      L@      �?       @      G@      @     �f@      "@     @V@      5@      �?      �?       @      $@                              @      "@      @      @       @                      ?@     �P@      �?      �?     �A@      @     �^@      *@     �_@      3@       @              4@     �E@                      $@             @X@      "@     �R@       @                      &@      7@      �?      �?      9@      @      9@      @     �I@      &@       @              4@     �E@      �?       @      D@             �`@      ,@     �K@      .@                      ,@     �A@      �?      @      :@              I@      *@      ;@      $@                      @      (@      �?       @      0@              ;@      @      *@      @                      @      7@              @      $@              7@      "@      ,@      @                      @       @              @      ,@             �T@      �?      <@      @                      @      @              @      "@             �E@              .@      @                              @                      @              D@      �?      *@      �?              1@     �l@      w@      <@      A@     �t@      N@     ��@     �g@     (�@     �q@      7@      @     �N@     �c@       @      @     �_@      1@     �t@      Q@     �p@     �]@      @      �?       @      3@                      1@              *@       @      (@      .@              �?              ,@                      $@              @      @      @      ,@                       @      @                      @              @      �?       @      �?               @     �M@      a@       @      @     �[@      1@     �s@      N@     �o@     �Y@      @       @     �J@     @V@      @      @     @T@      .@     �c@      M@     �_@      S@      @              @      H@      @      @      =@       @      d@       @     �_@      ;@              ,@     �d@     �j@      4@      ;@      j@     �E@     �m@      ^@     �q@      e@      1@      @      Z@     `b@      ,@      6@      b@      4@     �d@     �Q@     `g@      S@       @             �H@     �A@      @      &@      C@      @      H@      9@     �F@      ;@      �?      @     �K@      \@      &@      &@     �Z@      ,@     @]@      G@     �a@     �H@      @      &@     �O@     @P@      @      @      P@      7@     �Q@     �H@      X@      W@      "@      &@     �B@      G@      @      @      >@      3@      >@     �@@      C@      R@      "@              :@      3@               @      A@      @     �D@      0@      M@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ0�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�m�{TF@�	           ��@       	                    @����@�           ��@                           �?.�5Xh@�           0�@                           �?3����@)           `~@������������������������       �����1@q            �g@������������������������       �]��΍�@�            �r@                          �;@�<��@r             h@������������������������       ���KS9&@j            �e@������������������������       ��ӿ� @             2@
                           �?���Hx}@�            �w@                           @���H֢�?P             a@������������������������       ��Gr����?1            �S@������������������������       �d=Z�Cx�?            �L@                           @ќ�	a@�            �n@������������������������       ���Lz�@t            �f@������������������������       �*Ż�@/            �P@                           @�QM�-Z@�           H�@                           �?녬}��@�           ��@                            @�*(��;	@�           �@������������������������       ���{Q.	@%           �|@������������������������       ��R���(	@�           ��@                            @0�I��@	            z@������������������������       �
��g�@�            �o@������������������������       ����ߌ8@g            @d@                           �?�xB��@@$           �@                          �4@��Ơ��@�           (�@������������������������       ��p�N�@�            �v@������������������������       �ȧ
@@�            �s@                           @aYz�B@�           ��@������������������������       ����{v@           �z@������������������������       �v�~��.@t            @f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     0q@     `�@      =@      K@     �{@     �W@     ��@     `n@     ��@     �v@      0@      @     �R@     �a@      @      .@     @_@      4@     �s@     �S@      f@     �X@       @      @      N@      [@      @      ,@     �Z@      *@      ^@     @Q@      Z@     �Q@       @      @     �I@     �P@      @       @     �S@      &@      S@      M@     @Q@      L@      @      @      1@      ?@               @      A@      @      <@      @@      5@      0@       @              A@     �A@      @      @     �F@      @      H@      :@      H@      D@      @              "@      E@              @      ;@       @      F@      &@     �A@      ,@       @              "@      D@              @      5@       @      F@      &@      =@      (@                               @                      @                              @       @       @              .@      @@              �?      3@      @     �h@      $@     @R@      <@                              "@                      @       @     �W@      �?      .@      $@                               @                                     �L@              @      @                              �?                      @       @      C@      �?       @      @                      .@      7@              �?      .@      @     �Y@      "@      M@      2@                       @      4@                      $@             @U@      @     �C@      *@                      @      @              �?      @      @      2@      @      3@      @              8@      i@      z@      :@     �C@      t@     �R@     (�@     �d@      �@     �p@       @      6@     �a@     `m@      3@      >@     �k@     �H@     �q@      `@     �n@     �g@      @      6@      \@     @g@      1@      9@     �d@     �B@      g@     �U@      c@     �c@      @       @      G@     @P@       @      $@     @P@      3@     �O@      =@      Q@      T@              ,@     �P@     @^@      "@      .@     �Y@      2@     �^@      M@      U@     @S@      @              >@     �H@       @      @      K@      (@      X@     �D@     @W@      A@                      6@      9@      �?      @     �E@       @     �F@      :@     �P@      .@                       @      8@      �?       @      &@      @     �I@      .@      ;@      3@               @      M@     �f@      @      "@     �X@      9@     �|@      B@     �t@     @R@       @       @      <@     @Y@      @      "@     �F@      "@     �p@      ,@     �c@      D@       @              (@      L@      @       @      *@      �?     `f@      @     �S@      .@               @      0@     �F@      �?      @      @@       @     �U@       @      T@      9@       @              >@      T@      @              K@      0@     `h@      6@     �e@     �@@                      0@     �J@                     �@@      @     �c@      &@     �`@      1@                      ,@      ;@      @              5@      "@     �B@      &@      D@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�9lhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @*�n8P@�	           ��@       	                    �?Ӫ�I�@�           ȥ@                           �?>ҁ�V�@K           ��@                           �?�;2�)@�            �s@������������������������       �!I��=7@N            �`@������������������������       �~��[�@i            �f@                           @��|<�^@�           ��@������������������������       �p�у�;@0           �@������������������������       ��h(��@d            �c@
                          �5@a"5�]�@�           @�@                           @'7�}�C@�           ��@������������������������       ��'�S@�           �@������������������������       �\�(���@�            �w@                           �?��~�]	@           ؈@������������������������       ��P��߽	@%             O@������������������������       �&X]��@�           �@                          �2@�$�n�@�           ��@                           �?ڷɲw�@�            pq@                           �?z�Ԛ�=@G            @Y@������������������������       �2vsJ��@$             I@������������������������       ���k^ �?#            �I@                           @+b�]�@m            @f@������������������������       ��� !�@8             T@������������������������       ��4Ӯ�@5            �X@                           �?ʀn���@           p�@                          �8@<�>m!T@�            �j@������������������������       ��$�

@W             `@������������������������       �5ڐ�z@0            �T@                           �?4�&U�	@�           Ѓ@������������������������       ����Rn	@�            @o@������������������������       ���o��@�             x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@      �@      :@      M@      |@     �U@     ��@     �i@     P�@     �u@     �C@      $@     �j@     `x@      ,@     �B@     `s@      P@      �@     �a@      �@     @m@      :@      �?     �O@     �b@      @      @     �T@      (@     0v@      5@     `j@      Q@      @      �?     �@@     �O@      �?      @      D@      @      K@      ,@     �P@     �A@      @      �?      .@      7@      �?      @      0@      @      <@      $@      7@      $@      �?              2@      D@                      8@              :@      @     �E@      9@      @              >@      V@       @      @     �E@      "@     �r@      @      b@     �@@       @              8@      O@                      >@      "@     `o@      @      Z@      4@      �?              @      :@       @      @      *@              I@      @     �D@      *@      �?      "@     �b@     �m@      &@      ?@     `l@      J@     z@     @^@     �v@     �d@      4@              M@     �`@      @      ,@     �[@      3@     �q@     �K@     �n@     �U@      @             �@@     �S@      @       @     @U@      1@     `c@      @@     �d@     �N@      �?              9@      L@      �?      @      9@       @     @_@      7@     �T@      9@      @      "@      W@     @Z@      @      1@     @]@     �@@      a@     �P@     �]@      T@      *@      @      "@      @              @      (@      �?      @      @      $@      @      @      @     �T@     �Y@      @      &@     @Z@      @@     �`@     �N@     @[@     @S@      $@      @      Y@     �c@      (@      5@     �a@      6@     @n@      P@     @m@     @\@      *@      �?      .@      B@       @      @      ?@      �?     �W@      $@     �O@      5@              �?      �?      *@       @              (@      �?     �A@              ;@      "@              �?              @       @              (@      �?      &@              &@      @                      �?       @                                      8@              0@       @                      ,@      7@              @      3@              N@      $@      B@      (@                      @       @              �?      @              A@      @      2@      �?                       @      .@              @      *@              :@      @      2@      &@              @     @U@     �^@      $@      1@     @[@      5@     `b@      K@     `e@      W@      *@              3@      ;@              @      9@             �G@      ,@     �I@      6@                       @      4@              �?       @              B@      @     �C@      (@                      &@      @              @      1@              &@      "@      (@      $@              @     �P@     �W@      $@      $@      U@      5@      Y@      D@      ^@     �Q@      *@      @     �@@      B@      @      @      8@      "@      ?@      (@      I@     �A@      @      �?     �@@     �M@      @      @      N@      (@     @Q@      <@     �Q@     �A@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�,�Y^k@�	           ��@       	                   �:@�����L	@           ��@                          �6@6�[���@F           ܔ@                           �?cR���@?           ��@������������������������       ���wG@�            Pu@������������������������       ��i���u@o           �@                          �7@2!����@           z@������������������������       �)S5��@M            �^@������������������������       �G&��/	@�            pr@
                           @�T�
@�            �t@                           �? "���	@�             r@������������������������       �$l���@G            �[@������������������������       ���r1@	@l             f@                           �?�qXt}�@             D@������������������������       �      �?              @������������������������       �1�0�@             @@                           @�
GI�!@�           ��@                           �?�kK���@�           P�@                           �?��'�@q            �g@������������������������       ����Q?�@3            �V@������������������������       �5p���@>            �X@                           �?�/�x��@           �z@������������������������       ���@             @@������������������������       �B�� @�            �x@                           @t?D\@@(           ��@                           @��R��@�           x�@������������������������       ��&�G�@�           �@������������������������       ����J@!           �{@                           �?�VBiaR@I           �@������������������������       ��{[�@�             h@������������������������       �2!X/�Z@�            t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     �q@     ؀@      B@     �O@     �~@     �Q@     P�@      m@     Ј@     �u@      9@      ;@      d@     �j@      4@     �D@      q@      F@     Pp@     �a@     @p@      i@      4@      .@     ``@      f@      *@      ?@     �k@      >@      l@     �[@     `l@     �`@      1@      .@     @T@     �]@      @      5@      a@      .@     �f@     �R@      d@     @Y@      "@      @     �@@      K@      @      @     �J@      "@     �R@      =@     �A@      D@      �?      &@      H@      P@       @      2@      U@      @     @Z@     �F@     @_@     �N@       @              I@     �M@      @      $@     �U@      .@     �F@     �B@     �P@      A@       @              6@      *@      �?      @      =@      �?      @      @      8@      1@      �?              <@      G@      @      @     �L@      ,@     �D@      ?@     �E@      1@      @      (@      >@      C@      @      $@     �I@      ,@      B@      =@     �@@     @P@      @      @      <@     �@@      @      $@      H@      ,@      ?@      3@      ?@      N@      �?      �?      @      ,@      @      @      :@      &@       @      @      (@      :@              @      7@      3@      @      @      6@      @      =@      ,@      3@      A@      �?      @       @      @                      @              @      $@       @      @       @                      �?                                              @      �?       @              @       @      @                      @              @      @      �?      @       @      �?     �^@     @t@      0@      6@      k@      ;@     (�@     @W@     ��@     �b@      @              E@      W@      @      "@      R@      &@      d@     �F@     �^@      L@       @              0@      ,@              �?      4@      �?     �Q@      @     �H@      &@      �?              (@      "@              �?      (@              @@      @      0@      @                      @      @                       @      �?     �C@       @     �@@      @      �?              :@     �S@      @       @      J@      $@     �V@      D@     �R@     �F@      �?              @      @              @      @      �?      �?      @      �?      @                      7@     @R@      @       @     �H@      "@     @V@     �A@     @R@      C@      �?      �?      T@      m@      &@      *@      b@      0@      �@      H@     �y@      W@      @      �?     �I@     �c@       @       @     �V@      "@      {@      <@     Pr@      I@       @      �?      5@     �R@              �?     �G@       @     �s@      0@     �d@      ;@                      >@     �T@       @      �?     �E@      �?      ^@      (@      `@      7@       @              =@      S@      "@      &@     �K@      @     @b@      4@     �]@      E@      �?              @      A@      �?       @      .@      �?      S@      @      E@       @      �?              6@      E@       @      "@      D@      @     �Q@      ,@      S@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ3	$khG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@q*��kd@�	           ��@       	                    �?ɯ���@l           �@                          �3@�b��~{@�           x�@                          �2@rv[E^�@_           ��@������������������������       �md,@G� @           �z@������������������������       ���}��A@G            �[@                          �4@���Ծ@�             k@������������������������       ��&a�@@?            �W@������������������������       �ꔇA�@O            �^@
                           @d��Z�@           �@                           @�m[@�           ��@������������������������       ��iUol�@a            �b@������������������������       ��F��5@e           �@                           @ֹ0/�@�           x�@������������������������       �PjG=�@H           H�@������������������������       �{�oR@q            �d@                           @�,���@I           P�@                           �?q�*A��@�           p�@                           �?��v�_$@*           0}@������������������������       �/��Bh�@�             l@������������������������       �(�o:@�            @n@                           �?o^�[4	@�           $�@������������������������       �[�K}�8@�            �x@������������������������       �
�6t�{	@�           ��@                           �?�3Ъ�	@u             g@                            @��A
@6            �T@������������������������       �M���@&            �L@������������������������       �caa&<�@             9@                           �?���%]�@?            �Y@������������������������       �8�k8@            �D@������������������������       ���tn4@)            �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     Ѐ@      @@      J@      ~@     �S@     ��@      j@     (�@     �v@     �C@      @     @^@     �q@       @      6@     �m@      9@     ��@      W@     0}@     �d@      ,@              B@     �V@              @      M@      @     �u@      0@     `c@     �C@      @              7@      I@               @      C@       @     p@      $@      ^@      @@                      4@     �C@               @      ?@      �?     �k@      @     �S@      7@                      @      &@                      @      �?     �A@      @     �D@      "@                      *@     �D@               @      4@      @     �U@      @     �A@      @      @              @      0@                      &@             �C@       @      .@      @      @              $@      9@               @      "@      @      H@      @      4@       @              @     @U@     �g@       @      2@     `f@      4@     �w@      S@     �s@     �_@      &@      @      I@     �Z@      @      .@     �\@      ,@     �a@     �P@      _@     �R@      @      @      @      &@      @      �?      ;@      �?      <@      1@     �@@      ,@       @       @     �E@     �W@      @      ,@      V@      *@     �\@      I@     �V@      N@      @             �A@      U@       @      @      P@      @      n@      "@     �g@      J@      @              8@     �N@              �?     �F@      @     @i@      @     �a@     �A@      @              &@      7@       @       @      3@      @      C@      @     �G@      1@      �?      *@     @h@     p@      8@      >@     `n@     �J@     r@     @]@      s@     �h@      9@      &@      d@     �k@      4@      >@     @k@     �G@     �p@     @X@     @r@      g@      .@      �?     �D@     @Q@      @      @      O@       @     �W@      9@     @\@     �D@       @      �?      :@      C@       @      @     �@@      @      I@      &@     �B@      1@                      .@      ?@      @              =@      @     �F@      ,@      S@      8@       @      $@      ^@      c@      .@      9@     �c@     �C@     �e@      R@     `f@      b@      *@      �?     �C@      Q@       @      @      N@      "@     �I@      9@      P@     �P@       @      "@     @T@      U@      *@      5@      X@      >@     @^@     �G@     �\@     �S@      @       @     �@@      B@      @              9@      @      6@      4@      ,@      (@      $@       @      $@      (@      @              .@      @      @      $@      @      @      "@      �?      @      @      @              *@      @      �?      "@      @       @      "@      �?      @       @                       @              @      �?               @                      7@      8@      �?              $@      �?      .@      $@      "@       @      �?              $@      @                      @               @      @      @              �?              *@      1@      �?              @      �?      @      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJRV�1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �1@Ԉ�PV@�	           ��@       	                    @f��P	�@�           8�@                            @:Y�7��@�            0q@                            �?^�ƃ�@i             f@������������������������       �C�x���@Y            �b@������������������������       ��B�A� @             =@                           @�Y�@A            �X@������������������������       ����>(�@0             Q@������������������������       ���S!��@             >@
                           @����ơ�?�            @u@                           @	�ɕ��?�            �p@������������������������       �RѪ�O�?n            `d@������������������������       �މ2"8� @B            �Z@                            �?��,��?/            �Q@������������������������       ��+�[�.�?              H@������������������������       ��=Ú�6�?             7@                           @���0��@2           ĩ@                           �?�>S5	@�           <�@                            �?ۼ��QX	@�           ��@������������������������       ��P����@�             v@������������������������       �5�2�A	@�            pu@                          �:@����	@           `�@������������������������       �}=1�F�@q           ��@������������������������       ��Ξ��V	@�            0p@                          �7@�k��yw@b           L�@                           @��%�w�@k           ��@������������������������       ���,�@�            `l@������������������������       ���5��@�           h�@                          �<@���K�@�            0x@������������������������       �_LY��4@�            pr@������������������������       �������@@             W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@      s@     Ѐ@      @@     �F@     p}@      S@     ��@     �i@     p�@      x@     �A@              :@     @S@      �?       @     �D@              p@      =@     �b@     �@@      �?              4@     �C@      �?              4@             �T@      :@      P@      7@                       @      8@                      0@             �M@      ,@     �D@      .@                      @      5@                      "@              G@      &@     �C@      .@                      �?      @                      @              *@      @       @                              (@      .@      �?              @              7@      (@      7@       @                      @      (@      �?              @              5@      @      2@      �?                      @      @                      �?               @      @      @      @                      @      C@               @      5@             �e@      @     @U@      $@      �?              @      >@                      4@             @`@      �?      R@      "@      �?              @      ,@                      "@              Y@      �?      >@      @      �?               @      0@                      &@              >@              E@      @                               @               @      �?              F@       @      *@      �?                              �?               @      �?              @@       @      "@      �?                              @                                      (@              @                      5@     �q@     �|@      ?@     �E@     �z@      S@     ��@     @f@     Ȅ@     v@      A@      5@     �k@     �q@      7@      B@     0r@      M@      q@     `b@     s@     `n@      =@      @     �R@      X@      ,@      "@      \@      >@      ]@     �H@     �W@     �T@      $@      �?      D@      M@      @      @     �G@      *@     �O@      @@     �H@     �@@       @      @     �A@      C@      &@      @     @P@      1@     �J@      1@     �F@      I@       @      ,@     @b@     �g@      "@      ;@     `f@      <@     �c@     �X@     `j@      d@      3@      @      Z@     �d@      @      9@     �a@      4@      `@     �R@     `f@     @]@      0@       @      E@      9@      @       @     �C@       @      >@      7@      @@     �E@      @             �M@     �e@       @      @     `a@      2@     @|@      ?@     �v@     �[@      @              D@     ``@      @      @     �R@      *@     v@      $@     �p@     �Q@      @              *@      F@       @              ,@      $@     �Q@       @     �J@      0@       @              ;@     �U@      @      @      N@      @     �q@       @     �j@     �K@       @              3@     �E@      �?       @     @P@      @     �X@      5@      W@     �C@      �?              &@      :@      �?       @      G@      @     �U@      3@     @S@      6@      �?               @      1@                      3@      �?      *@       @      .@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ǩhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�ȮyT@�	           ��@       	                    �?`M����@�           |�@                           �?�-�᥆@!            �@                            �?��k�ۇ@�            pq@������������������������       ��|lnޕ@S             _@������������������������       ����t�@X            `c@                          �8@�r$m�8@v           H�@������������������������       �h�h�]C@B            @������������������������       ��%���@4            �U@
                           @�[S�ߺ@�           x�@                           @�_8�|@           ��@������������������������       ��.�V@�            �t@������������������������       �*��-t$@C           ��@                          �5@}휌$.@�            �m@������������������������       ����`�@A            �V@������������������������       �*�IS@]            �b@                           @2�h�� @�           ,�@                           �?!�����@(           ȋ@                           �?�[L��@�            `n@������������������������       ��ч�9@S            �^@������������������������       ��_�@D             ^@                           �?J0�"W	@�           0�@������������������������       ��s� �8	@%             Q@������������������������       ����$	@l           �@                           @bi1E�5@�             q@                           @�}�)Ĺ@S             a@������������������������       ��n:���?            �E@������������������������       �
�e�@<            �W@                           @*/�]�@X             a@������������������������       ��]�˪��?1            �R@������������������������       ���~�F�@'            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     Pr@     x�@      @@      L@     �|@     @S@     H�@     @m@     �@     `w@      =@      @     `i@     �v@      &@      E@     Ps@     �I@     �@     `f@      �@     `n@      5@      @      K@     �Z@       @      @     �S@      @      u@     �B@     @f@      J@      @      @      ;@      H@      �?      @      A@      �?      N@      3@      I@      =@       @      @      @      @@              �?      &@      �?      9@      @      ?@       @                      4@      0@      �?      @      7@             �A@      ,@      3@      5@       @              ;@     �M@      �?      �?      F@      @     @q@      2@      `@      7@      @              :@     �H@      �?      �?     �C@       @     �o@      *@     �Y@      (@      �?              �?      $@                      @      @      8@      @      :@      &@       @      @     �b@     @p@      "@      B@     �l@     �F@      {@     �a@      w@     �g@      0@      @     @\@     �m@       @      A@      i@      B@     @x@     @Z@      u@     `e@      *@      �?      ?@      @@       @      *@     �G@      $@      N@      <@      R@      B@      �?       @     �T@     �i@      @      5@     @c@      :@     �t@     @S@     �p@     �`@      (@              B@      7@      �?       @      >@      "@      G@     �B@      @@      4@      @              "@      "@               @      $@      @      :@      @      &@      *@       @              ;@      ,@      �?              4@      @      4@     �@@      5@      @      �?      ,@     �V@      d@      5@      ,@     �b@      :@      q@     �K@     �k@     ``@       @      ,@     �S@      a@      1@      *@     �^@      8@     �e@      I@     �`@     �]@      @              ,@      D@       @      @      A@      �?     @S@      .@      B@      3@                      @      4@       @      @      ,@      �?     �C@       @      5@      "@                      "@      4@              �?      4@              C@      @      .@      $@              ,@      P@      X@      .@       @     @V@      7@     �X@     �A@     @X@      Y@      @      @      *@      "@              �?      (@       @      @      @      "@      @       @      "@     �I@     �U@      .@      @     @S@      5@     �W@      =@      V@     �W@      @              (@      8@      @      �?      <@       @     @X@      @      V@      (@      �?               @      &@              �?      "@       @     �O@      @      B@       @                       @      @                               @      3@              *@                              @      @              �?      "@              F@      @      7@       @                      @      *@      @              3@              A@              J@      $@      �?               @      @                       @              6@              B@       @      �?               @      $@      @              &@              (@              0@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Ӣ~�*@�	           ��@       	                     @��	�ک@H           ��@                           �?Z����]@:           L�@                          �<@����s�@           pz@������������������������       ��3%�mH@�            �w@������������������������       ��	<��C@             F@                          �2@eFI���@2           `�@������������������������       �-��X�*@i             e@������������������������       �=���A	@�            �@
                           �?�#���@            �@                          �<@�j	���@�            �k@������������������������       ������O@z            �h@������������������������       ��%"�Kq@             7@                           �?X�սͤ	@�           @�@������������������������       ���K�a@$             K@������������������������       �[����U	@b           ��@                          �4@�w�<U@p           ț@                          �1@�޷ �@b           ��@                           @�z�H%��?�            0w@������������������������       ���I�u��?�            �r@������������������������       ���'D���?,            @Q@                           @^ܷ2��@x           �@������������������������       ���)��e@`            �a@������������������������       �4��a�@            {@                          �7@��a�p5@           ��@                           @����q�@�            �x@������������������������       ��Җld@�            �q@������������������������       �i�v�J@B            �Z@                           @0�W	u�@           `{@������������������������       ��&�P/@�             n@������������������������       ���#�@t            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        "@      r@     8�@      @@     �J@     �{@     @W@     |�@     �j@     H�@     �v@      =@      "@     �i@     Ps@      :@     �B@     �r@      P@     0x@      e@     `w@      m@      6@      �?      `@     �d@      "@      2@      g@      G@      m@      ]@      m@     @c@      &@      �?     �F@     �G@      �?      �?     �J@       @      [@      2@     �Y@      D@      @      �?     �B@      F@      �?      �?      H@       @      [@      1@      X@      7@      �?               @      @                      @                      �?      @      1@      @             �T@     �]@       @      1@     �`@      F@      _@     �X@     @`@     �\@      @              "@      5@                      9@      �?     �G@      .@     �B@      *@                     �R@     �X@       @      1@     �Z@     �E@     @S@     �T@     @W@     @Y@      @       @     �S@     �a@      1@      3@     �\@      2@     `c@      J@     �a@     �S@      &@              2@      A@              @     �A@             @Q@       @      E@      $@                      2@      ?@               @      ;@             �O@      @      E@      @                              @               @       @              @      �?              @               @      N@     @[@      1@      .@      T@      2@     �U@      F@     �X@     @Q@      &@      @      @      &@              �?      "@      �?              *@      @      @       @      @      K@     �X@      1@      ,@     �Q@      1@     �U@      ?@     �W@     �P@      "@              U@     @n@      @      0@     `b@      =@     ��@     �F@     0y@     ``@      @              D@      ^@       @       @     �D@      @     �{@      2@     �i@      M@      �?              "@     �F@              @      ,@             �h@       @     �S@      3@      �?              "@     �A@                      ,@              d@              Q@      ,@      �?                      $@              @                     �B@       @      &@      @                      ?@     �R@       @      @      ;@      @      o@      0@      `@     �C@                      4@      ?@                      @      @      F@      @      ;@      @                      &@      F@       @      @      6@       @     �i@      $@     @Y@     �@@                      F@     �^@      @       @     �Z@      7@     �k@      ;@     �h@     @R@      @              0@     �Q@      �?       @     �H@      .@      _@      @      U@      7@      @              @      J@                      ?@      ,@     �X@       @      Q@      ,@                      "@      2@      �?       @      2@      �?      :@      �?      0@      "@      @              <@      J@      @      @     �L@       @     @X@      8@      \@      I@      �?              0@      ?@                      @@      @     �O@      "@     �O@      6@      �?              (@      5@      @      @      9@      @      A@      .@     �H@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ[TIhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�a�3�r@�	           ��@       	                   �2@�= ��@{           �@                          �1@f�wU$R@H           0�@                           �?��v1@�            �r@������������������������       �lg�i7b@L             ^@������������������������       ���hsC@t            �f@                            @D��|pU@�             k@������������������������       �ܩr��@I            @\@������������������������       �[�.�@?            �Y@
                          �;@Ӳ�l	@3           $�@                           �?��1�8	@x           ؕ@������������������������       �R��e��@           �z@������������������������       �:"���	@e           8�@                           @�QB���	@�            0q@������������������������       �D�FHm	@            �h@������������������������       ���:�1@<            �S@                           �?TDG�q)@.           �@                          �5@�Gk�S� @s           ��@                           @`Ej���?
           �y@������������������������       ���ܼ���?�            �q@������������������������       �Ҽ���O@R            �_@                           @	%bq@i            �d@������������������������       � 2��5@�?9             W@������������������������       �T����@0            @R@                           �? �ٲn@�           �@                           @�P}'@S           `�@������������������������       �냪��+@�             v@������������������������       �*�׋�f@~            @i@                           @pH[1�a@h           ��@������������������������       �g4� ��@V           @�@������������������������       ��R
Ԋ�@             D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     0s@     `�@      ?@     �O@     �|@     @U@      �@     �k@     ��@     �w@      ;@      2@     �i@     �s@      0@      H@     �s@     �R@     pw@      g@     �u@     �p@      6@       @     �B@     �Q@      �?      @      P@      @      b@     �B@     @Y@      J@              �?      6@     �D@      �?      �?      @@      �?      X@      2@     �P@      7@              �?      @      4@      �?              1@      �?      E@       @      *@      &@                      0@      5@              �?      .@              K@      $@     �J@      (@              �?      .@      =@              @      @@      @      H@      3@     �A@      =@                      @      $@                      .@       @      ?@      0@      3@      ,@              �?      "@      3@              @      1@      @      1@      @      0@      .@              0@      e@     �n@      .@      F@     `o@     @Q@     �l@     �b@      o@      k@      6@      @     �`@      j@      .@      >@     @k@      J@     �i@     @^@     `l@     �c@      3@             �H@      N@       @       @      L@      @      W@      8@     @Y@      @@       @      @     �U@     �b@      *@      6@     @d@     �G@     �\@     @X@     �_@     �_@      1@      "@     �@@     �A@              ,@     �@@      1@      8@      ;@      5@     �M@      @      "@      8@      @@              $@      2@       @      1@      0@      ,@     �F@      @              "@      @              @      .@      "@      @      &@      @      ,@               @     �Y@     @j@      .@      .@     �a@      $@     h�@     �B@      |@     @\@      @              4@     �P@       @      �?      ?@      @     �q@      @     �a@      .@       @              0@      I@              �?      0@             �k@      @     �V@       @       @              "@      A@                      "@             `e@              K@      @                      @      0@              �?      @             �I@      @     �B@      @       @              @      0@       @              .@      @      P@      @     �I@      @                      @       @                      @      �?     �E@              =@       @                      �?       @       @              "@       @      5@      @      6@      @               @     �T@      b@      *@      ,@     �[@      @     �t@      ?@     @s@     �X@      @       @      E@      S@      @      &@      M@             @c@      *@      d@     �@@       @       @      4@     �K@      @      @     �C@             @T@      @      _@      5@                      6@      5@               @      3@             @R@      "@      B@      (@       @              D@      Q@       @      @     �J@      @     �f@      2@     �b@     @P@      �?              =@      P@      @      @     �G@      @      f@      0@     �a@     �O@      �?              &@      @      @              @      @      @       @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ	�z	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�?��0@�	           ��@       	                    �?�ٻ�@�           �@                           �?w��3@/            �@                            �?�ٌC{d@w            �h@������������������������       �f���ԝ@(             P@������������������������       ���0��@O            �`@                            �?�˝�w�@�            �s@������������������������       ���.��@X             b@������������������������       ���n��U@`            �e@
                          �8@xF@��@�           �@                          �1@�̸�57@�           (�@������������������������       ��,6TX�?y            �g@������������������������       �%i���F@           pz@                           @@��e��@D             W@������������������������       �����K@<            �T@������������������������       �=��,@             $@                           �?��(��@�           �@                           @S��@}             i@                          �5@c^N9u<@]            �b@������������������������       �{�ℙ@$             M@������������������������       ����Pm&@9            @W@                          �6@���f�@             �H@������������������������       �B�P$@            �A@������������������������       �騼����?             ,@                            �?,_:u�@8           ��@                          �3@�o��A�@�           ؄@������������������������       ����� @�            `j@������������������������       ��ِQ\�@&           �|@                           @���u�@�           ��@������������������������       �G�ʏ~�@g           ԛ@������������������������       ��t�rP@!             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     @s@     p�@      6@      I@     �~@     @P@     ��@     �k@     ��@     `v@     �A@       @     �T@     @d@              (@      ^@       @     0{@     �J@      p@     �S@      @       @      K@      U@               @     �P@       @      [@     �A@     �V@      M@      @       @      *@     �C@                      4@              L@       @      C@      2@       @       @       @      (@                      @              4@      �?      0@      @       @              &@      ;@                      .@              B@      @      6@      ,@                     �D@     �F@               @     �G@       @      J@      ;@      J@      D@       @              .@      5@              @      7@              6@      .@      4@      7@       @              :@      8@              @      8@       @      >@      (@      @@      1@                      =@     �S@              @     �J@      @     pt@      2@      e@      5@      �?              <@     @Q@              @      G@       @     �r@      ,@     @a@      ,@                       @      1@               @      "@             �[@      �?      F@      @                      :@      J@               @     �B@       @     `g@      *@     �W@      $@                      �?      "@                      @      @      =@      @      >@      @      �?                      "@                      @      @      <@      @      =@      @      �?              �?                              �?      �?      �?      �?      �?      @              &@      l@     �z@      6@      C@      w@     �L@     ��@      e@     x�@     pq@      >@      �?     �@@      2@              @      D@      @      "@      5@     �C@      8@      @      �?      @@      0@              @      ?@      @      @      0@      .@      5@      @              @       @              @      (@       @      �?      @       @      *@              �?      <@       @              �?      3@       @      @      &@      @       @      @              �?       @                      "@      �?      @      @      8@      @                               @                      "@      �?      @       @      0@      �?                      �?                                                      @       @       @              $@      h@     �y@      6@      @@     �t@      J@     ��@     �b@     �~@     �o@      :@      �?     �I@     @V@       @      *@     @U@      3@     `e@      M@     �[@      O@      @               @      5@              �?      8@       @     �T@      @      E@      6@      �?      �?     �E@      Q@       @      (@     �N@      1@      V@     �I@     @Q@      D@      @      "@     �a@     t@      4@      3@     `n@     �@@     �v@     �V@     �w@      h@      5@       @     @`@      t@      4@      3@     �l@      @@     @v@      V@     w@     �g@      4@      �?      &@      �?                      (@      �?      @       @       @      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJA�#chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?:��.-@�	           ��@       	                   �4@�E*�hc@�           ��@                           @�V��y@�           x�@                           �?��(o@�            0s@������������������������       �Nރ޺@|             k@������������������������       �#C]��@=            �V@                            �?�v�%��?�            �u@������������������������       ��d��� @n             g@������������������������       �Y�j��?j            �d@
                           �?� ��@a           ��@                          �6@?��I@�            �o@������������������������       �T�m��B@5             R@������������������������       �X��a�@t            �f@                           @_n���.@�            pq@������������������������       �V����@;            �W@������������������������       �b�u)�/@}             g@                            @Haj@�           H�@                           @Sn���@�           0�@                          �2@u����L	@`           �@������������������������       ��Go�g8@u            `f@������������������������       �h�	A	@�           p�@                           @UkKT��@^           X�@������������������������       �텓�l@s            `g@������������������������       ��eN61P@�           ��@                           �?��lbQ�@�           ��@                           �?����1�@�            �s@������������������������       ��@3=gZ	@q            `g@������������������������       �ۧߜ��@T            �`@                           @�R�Ǎ@)           �}@������������������������       ���$�p @F            @Z@������������������������       �%��]�r@�             w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     �s@     ��@      =@      M@     @|@     �R@     ��@     �j@     8�@      v@      ;@      �?     @U@     `e@      @      @     �W@       @     �y@     �@@     �q@      V@       @              B@     �S@              @     �C@      �?     �q@      .@     �c@     �F@      �?              5@      D@              �?      <@      �?     �W@      $@     �S@      A@                      ,@     �B@                      3@      �?     �O@       @     �F@      =@                      @      @              �?      "@              ?@       @     �@@      @                      .@      C@               @      &@             `g@      @     �S@      &@      �?              *@      7@               @      @             �V@      �?     �C@      $@                       @      .@                      @              X@      @     �C@      �?      �?      �?     �H@     @W@      @      @      L@      @     ``@      2@      `@     �E@      �?      �?     �B@      G@      @      @     �C@      �?      C@       @     �F@      @@      �?              1@      @       @              @              1@      @      0@      @              �?      4@     �C@      �?      @     �A@      �?      5@      @      =@      :@      �?              (@     �G@                      1@      @     @W@      $@     �T@      &@                       @      @                       @      �?      ;@      @      @@      @                      @      D@                      "@      @     �P@      @     �I@      @              "@      m@     px@      :@     �I@     Pv@     �P@     ��@     �f@     X�@     �p@      9@      @     �c@     q@       @      B@     @o@     �H@     �{@     �`@     @x@      f@      0@      @      W@     �^@      @      9@     �c@      D@     @_@     �Y@     �`@     �Z@      (@      �?      0@      1@                      :@      �?     �K@      6@      8@      .@       @      @      S@     @Z@      @      9@     @`@     �C@     �Q@     @T@     �[@      W@      $@             @P@     �b@      �?      &@     �W@      "@     �s@      =@     �o@     �Q@      @              $@      <@      �?      @      (@      @      M@      (@     �D@      ,@                     �K@     �^@              @     �T@      @      p@      1@     �j@      L@      @      @     �R@     �]@      2@      .@     �Z@      2@     @_@     �H@     �d@     �U@      "@      �?      8@      B@      0@      &@     �F@      @     �I@      *@     �Q@      E@      @      �?      7@      4@      *@      $@     �B@       @      1@      @      <@      ;@      @              �?      0@      @      �?       @      @      A@      "@      E@      .@              @     �I@     �T@       @      @      O@      *@     �R@      B@     @X@     �F@      @      �?      *@      4@              �?      ,@      @      @      .@      6@      @      @       @      C@      O@       @      @      H@      @      Q@      5@     �R@     �D@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?U�j�@�	           ��@       	                    �?$����@            ē@                          �<@�Z|�[�@=           �@                          �1@Q���-@            |@������������������������       �r����(@1            �U@������������������������       �I�a��@�            �v@                            �?}���_@             �L@������������������������       ��>B֣@             ?@������������������������       �F�uz�@             :@
                          �3@��ʦ�&@�           ��@                            @�@����?�            �x@������������������������       �ͱ.Ȉ�?�            �t@������������������������       �Bl�K�?*             N@                           �?���}?�@�            �v@������������������������       �*O �n@�            @k@������������������������       ��u�z�@c            @b@                            @D��a�	@p           ��@                           @[����@�           p�@                           �?�+��B	@3           ��@������������������������       ���G���	@�           H�@������������������������       �*���/^@�            �r@                          �7@sl/��@\           @�@������������������������       �8�G��,@�           Ȇ@������������������������       �Z�V��@�            �m@                           �?ƿ�'�@�           ��@                          �8@bh����@+            �O@������������������������       �mM<'�j@            �D@������������������������       �H��/X�@             6@                           �?si��a@�           �@������������������������       ������	@           0{@������������������������       ��m��e�@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �q@     ��@      <@     �K@     @{@     �W@     ��@     �j@     ��@     `v@      2@              S@      d@       @      $@     �X@      "@     �}@      F@     �r@     @U@      @             �I@     �S@      �?      $@     �O@       @      _@      A@      Y@     �D@      @             �F@     �R@      �?      @      K@       @     @^@      >@     @V@      :@      @               @      &@                      1@             �A@      @      0@       @                     �E@     �O@      �?      @     �B@       @     �U@      :@     @R@      8@      @              @      @              @      "@              @      @      &@      .@                      @      @                                      �?       @      @      *@                                              @      "@               @       @      @       @                      9@     �T@      �?             �A@      @      v@      $@     �h@      F@      �?              &@      =@                      "@             �h@       @     �^@      6@      �?              $@      =@                      @             �d@       @     �X@      4@      �?              �?                               @              @@              7@       @                      ,@      K@      �?              :@      @     �c@       @      S@      6@                       @      >@                      1@      @     @\@      @      ?@      $@                      @      8@      �?              "@      @     �E@       @     �F@      (@              .@     �i@      w@      :@     �F@      u@     @U@     `�@     `e@     0�@     q@      ,@       @     �`@     �o@      *@      :@     �m@     �M@     �{@     �`@     @x@      g@      "@       @     �T@     �^@       @      2@     @a@     �G@     @^@     �Z@     �b@     �Z@       @       @      L@     �V@       @      (@     @W@      >@     �O@     �R@     �T@     �V@       @              :@     �@@              @     �F@      1@      M@      @@     �P@      .@                      J@      `@      @       @     �X@      (@      t@      :@     �m@     �S@      �?              D@     �Y@      @      @      M@      &@     0q@      ,@     �c@     �M@                      (@      :@              @      D@      �?     �F@      (@     �S@      4@      �?      @     @R@      ]@      *@      3@     �Y@      :@     `b@      C@     @`@      V@      @      �?      @      ,@              @      "@      @      �?      &@      @      @      @              @      $@              @      "@      @              @      @       @              �?      @      @                                      �?      @      @       @      @      @     �P@     �Y@      *@      0@     @W@      7@     @b@      ;@     �^@      U@       @      @      I@     �M@      (@      0@      R@      6@     �J@      3@     �N@     �O@       @              0@     �E@      �?              5@      �?     @W@       @      O@      5@        �t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ8�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?xS�mE@�	           ��@       	                    @�(e���@�           ��@                          �<@�A]��@�           8�@                           �?�۵i�$@r           h�@������������������������       ��3�v�@�             q@������������������������       ���HO�@�            �s@                           �?������@%             M@������������������������       �7M;ߜ@             @@������������������������       �b�ܵ@             :@
                          �4@֝t�G@a           �@                           �?n���?�            �s@������������������������       ��I s�.�?t            �e@������������������������       ��V
�d&�?`            �a@                            @.bN��E@�            �l@������������������������       �JHG:V@t            �g@������������������������       �������?             E@                           @�v��@�           B�@                          �:@&A��	@�           T�@                           �?�%~A��@           ��@������������������������       �����b	@2           �@������������������������       ��i̶�S@�            �u@                            �?���J�#
@�            Ps@������������������������       �AT}�8	@;             X@������������������������       ���	@�            �j@                           @��T8�x@�           0�@                          �<@x\�F7@�           ȑ@������������������������       �F�B�@�           ��@������������������������       ��m��f@*            �P@                           6@�c,��J@             :@������������������������       ��k�0��?             &@������������������������       �������@             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     ��@      B@      C@     �{@     �W@     �@     `j@     h�@     @w@      ;@      �?     �R@     �b@      @      "@     �Y@      *@     `z@      F@     pq@      V@      @      �?      N@     �S@      @      "@      S@      @     `d@     �A@     �b@      P@      @      �?     �K@      R@      @      @     �P@      @     `d@      8@     `a@     �I@       @      �?      <@      <@      @      @     �C@      @      V@      ,@      C@      8@      �?              ;@      F@              @      ;@       @     �R@      $@     @Y@      ;@      �?              @      @               @      $@                      &@      $@      *@      �?              @      @              �?       @                      @      @      "@                      �?       @              �?       @                      @      @      @      �?              ,@     @R@      �?              :@      @     0p@      "@     @`@      8@       @               @      A@                      &@             �f@      @      P@      $@       @              @      4@                      "@              Z@      @      =@      @                      @      ,@                       @             @S@       @     �A@      @       @              @     �C@      �?              .@      @     �S@      @     �P@      ,@                      @     �A@      �?              .@      @      I@      @      M@      ,@                       @      @                                      <@               @                      5@     `l@     �w@      @@      =@      u@     �T@     �@     �d@     ��@     �q@      6@      5@     �d@     @k@      :@      7@     @m@     �P@     �k@      b@     �m@     `f@      5@      @     �_@     �h@      4@      2@     �g@      I@      h@     �Z@     @j@     �]@      .@      @     @X@     `a@      2@      .@     @b@      A@     @]@     �S@     �a@     �V@      .@              =@     �L@       @      @     �E@      0@      S@      <@     �Q@      ;@              .@     �C@      6@      @      @     �F@      1@      <@      C@      ;@     �N@      @       @      @      @      �?      �?      2@      @      @      4@       @      0@      @      *@      A@      .@      @      @      ;@      $@      7@      2@      3@     �F@                      O@     @d@      @      @      Z@      .@      v@      6@     �t@     @Z@      �?              M@      d@      @      @     @Y@      "@      v@      4@     t@     �Y@      �?              H@     �b@      @      @      W@      "@     �u@      4@     0s@     �V@      �?              $@      $@       @              "@               @              ,@      *@                      @      �?                      @      @               @       @       @                                                              @                      @       @                      @      �?                      @       @               @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{�]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@sm�@�H@�	           ��@       	                    @k�b`�J@           ��@                           �?+�/�a@8           H�@                           �?���@�            @s@������������������������       �h��_?d@�             j@������������������������       �h𡧱@=            �X@                          �2@E��h8@y           ��@������������������������       �?AJ-�@�             p@������������������������       ���Kҙ�@�            Ps@
                            �?H3�}@G           �@                          �2@�*��BC@7           @}@������������������������       �@SK��@�             q@������������������������       ��~[@�            @h@                           @%ۓ�a@           �z@������������������������       �����Ȍ @�            �r@������������������������       ��u�%�@R            �_@                           @�Z��_@?           ��@                           �?ݚ�[X	@D           ��@                           �?f�Y�$@�             u@������������������������       �H��G@�             p@������������������������       ��'<u�@6             T@                            @K�����	@j           ��@������������������������       ���g�	@}           ��@������������������������       �B��8iy@�            �v@                           @����|@�           x�@                           �?�#�g:@^           ��@������������������������       ���ֈ��@�            @m@������������������������       �6��;�H@�            �t@                           @��3D@�            �o@������������������������       ��è�R@@�            �l@������������������������       �K�Rα@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     @�@      ,@     �P@      |@     @X@     (�@     �n@     h�@     �u@      <@      @      [@      k@      @      3@      d@      1@     X�@     �V@     0x@     �`@      $@      @     �O@      ^@      �?      $@      Z@      ,@     �i@     �R@     �e@     �W@       @              :@     �B@              �?      9@              Y@      9@     @Q@      8@      �?              2@      ;@              �?      0@              Q@      5@      B@      5@      �?               @      $@                      "@              @@      @     �@@      @              @     �B@     �T@      �?      "@     �S@      ,@     �Z@     �H@      Z@     �Q@      @       @      0@      G@              @      >@       @      M@      7@     �H@      ;@              @      5@     �B@      �?      @     �H@      (@      H@      :@     �K@      F@      @             �F@     @X@      @      "@      L@      @     �y@      0@     �j@     �C@       @              1@     �D@      �?      @      D@      �?     �i@      &@      ^@      =@                      (@      5@      �?      @      2@      �?      a@      @      L@      6@                      @      4@                      6@              Q@       @      P@      @                      <@      L@       @      @      0@       @      j@      @     �W@      $@       @              5@      D@              @      "@       @      d@       @     �L@      @       @              @      0@       @              @             �H@      @     �B@      @              "@     `f@     �t@      $@      H@      r@      T@     �w@     @c@     �z@      k@      2@      "@     �`@     `j@      "@      E@     �h@     �O@     `d@     �_@     �i@      c@      ,@      �?     �G@     �J@              @     �A@      @     �R@      .@     �Q@      9@      @      �?     �B@     �F@              @      >@      �?      H@      ,@     �I@      6@      @              $@       @                      @      @      ;@      �?      4@      @      �?       @     �U@     �c@      "@      B@     �d@     �L@      V@     �[@     �`@      `@      $@      @     �N@     �T@      @      8@      Y@      G@      M@     �T@     �T@     @R@       @       @      :@      S@      @      (@      P@      &@      >@      =@     �I@     �K@       @             �F@      _@      �?      @     �V@      1@     �j@      <@     �k@     �O@      @              5@     �U@      �?      @     @P@      ,@     @d@      (@      e@      =@                      @     �H@                      4@      @     �S@       @      Q@      "@                      1@     �B@      �?      @     �F@      &@     �T@      $@      Y@      4@                      8@      C@               @      :@      @     �J@      0@     �J@      A@      @              1@      B@               @      4@              J@      *@      I@      A@      @              @       @                      @      @      �?      @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�	 {>z@�	           ��@       	                    �?oN��@i           F�@                          �<@ODo2@�           ��@                            @k�I#�@o           8�@������������������������       �O��ґ�@�            pv@������������������������       �����(Q@�             l@                          �=@����@#            �K@������������������������       �x1���?             4@������������������������       ��=C�9{@            �A@
                          �5@sB��M�	@�           ��@                           �?�+�a@�           P�@������������������������       �'��T�@B           �~@������������������������       ���0(s@�             l@                           @ 	8��	@
           ؊@������������������������       ��W�
@J           ��@������������������������       �$C�7��@�            `t@                            �?=��N�+@7           ��@                          �5@ �F��@�            px@                           �?������?�            `o@������������������������       �6�YU��?6            �V@������������������������       ����D�@g             d@                          �7@.>�ǇY@U            �a@������������������������       ����`@             �J@������������������������       �M�Fo�@5            �U@                            @/��?@E           |�@                           @�iSTq@�           ��@������������������������       ���>.�@�           4�@������������������������       � �m�)�@             6@                           @W.��@�            �o@������������������������       �X�Uh��?T            �`@������������������������       ����V_@O            �]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     0r@     ؀@      A@      K@     p{@      X@     H�@     @n@     ��@     �w@     �B@      (@      j@     �t@      7@     �C@      s@     �Q@     v@      i@     pw@     `p@      =@              L@     �W@      �?      @     @Q@      $@     @c@      ;@     �c@      O@      @              J@     �U@      �?      �?     @P@      $@      c@      2@     �b@     �F@      @              B@      G@              �?     �D@      $@     �U@      *@     @X@      9@      @              0@     �D@      �?              8@             �P@      @     �I@      4@                      @      @               @      @              �?      "@      "@      1@       @                      @                                                      @      &@                      @      @               @      @              �?      "@      @      @       @      (@      c@     �m@      6@      B@     �m@     �N@     �h@     �e@     @k@      i@      8@      @     �B@      \@       @      ,@     @Z@      2@     �`@     �R@      `@     �R@      @      @      A@      P@      @      @     @T@      2@     �P@     �I@     �V@      N@      @              @      H@      @      @      8@             @P@      8@     �B@      ,@               @      ]@     �_@      ,@      6@     �`@     �E@     �P@     �X@     �V@     �_@      1@      @      U@     @P@      &@      .@     �V@      @@      A@     �I@      L@     �R@      .@      @      @@     �N@      @      @      E@      &@     �@@     �G@      A@     �I@       @             �T@     �i@      &@      .@     �`@      9@     @�@      E@     z@     �\@       @              3@      F@      @              9@      (@     �d@      &@     �U@      8@                      @      :@                      (@             �_@      @      P@      $@                               @                                      M@              6@      @                      @      2@                      (@             @Q@      @      E@      @                      (@      2@      @              *@      (@      C@      @      7@      ,@                       @      "@      @              @      �?      4@               @      @                      @      "@                      "@      &@      2@      @      5@      "@                     �O@     `d@      @      .@      [@      *@     0~@      ?@     �t@     �V@       @             �J@      b@      @       @     �W@      (@     �w@      :@     @p@     @R@      @             �G@      b@      @       @      V@      @     pw@      8@     @p@     �Q@      @              @                              @      @      �?       @               @                      $@      2@      �?      @      ,@      �?     �Z@      @     �Q@      1@       @              @      @                       @             �P@              F@       @       @              @      &@      �?      @      @      �?     �D@      @      :@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��B@�	           ��@       	                     �?S:R��n@�           ��@                           �?+�5D��@�           ��@                          �;@�.Q|�l@�            �o@������������������������       ��=��%C@�            �j@������������������������       �Ls�@�@             D@                          �8@�J��(@�            py@������������������������       �R�-]@@�             v@������������������������       ���I��@            �J@
                           �?.����@Z           Ѐ@                          �7@�E]�(@�            �i@������������������������       ���C��@c             c@������������������������       ��m�-r@'             K@                          �3@�/
�� @�            �t@������������������������       � ]QZ%<�?d            �d@������������������������       ����9#@l            �d@                           @�Q.��#@�           4�@                          �6@/"-b�|	@�           ��@                          �5@6�����@&           �@������������������������       �@��@�           �@������������������������       ���ɤ@X            �`@                          �:@� �/��	@�           ��@������������������������       �%�Z@�	@�            �w@������������������������       ��F7烺	@�            �q@                          �6@�I� ��@�           l�@                          �4@ �w1�@            �@������������������������       �X���L�@|           ��@������������������������       ��eeB6�@�            �i@                           @�]6��@�            pu@������������������������       ���S2#@�            �k@������������������������       ���WK�@S            �^@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     P�@      <@     �M@     p}@     @T@     `�@      i@     (�@     �w@     �A@      �?     �R@     �d@      @      @     �Y@      &@     �{@      A@     �p@      U@      @      �?     �D@     @W@      @      @      I@      $@      m@      ,@     �b@      M@       @      �?      9@      B@      @      @      :@       @     �L@      &@     �J@     �@@       @              5@      ?@      @       @      8@              K@      "@      I@      2@       @      �?      @      @              @       @       @      @       @      @      .@                      0@     �L@      �?              8@       @      f@      @     @X@      9@                      0@     �H@      �?              7@      @      d@      �?     �U@      ,@                               @                      �?      @      .@       @      &@      &@                     �@@      R@      �?       @      J@      �?     �i@      4@     @^@      :@      @              3@      D@      �?              A@      �?      E@      .@      B@      2@                      &@      >@                      4@      �?      @@      "@     �@@      0@                       @      $@      �?              ,@              $@      @      @       @                      ,@      @@               @      2@             �d@      @     @U@       @      @              @      "@                      @              Y@      @     �D@      �?      @              &@      7@               @      ,@             @P@              F@      @              *@      j@     Px@      7@      J@     w@     �Q@     ��@     �d@     ��@     �r@      >@      (@     @c@     �m@      3@     �E@     �n@      K@     �g@      a@     �l@     �g@      ;@      @     �T@     @^@       @      ;@     �`@      2@     @b@     �P@     �a@     �Z@      $@      @     �K@     @Z@      @      5@     @]@      0@      `@      N@     @`@      T@      $@      �?      <@      0@       @      @      1@       @      1@      @      *@      :@              @     �Q@     @]@      &@      0@      \@      B@     �E@     �Q@     @U@     �T@      1@              C@     �T@       @      @      P@      2@      :@     �A@     �M@      ?@      ,@      @     �@@     �A@      @      "@      H@      2@      1@      B@      :@     �I@      @      �?      K@     �b@      @      "@     �^@      0@     pw@      =@      s@      [@      @              A@      W@      @      @     @R@      &@     �r@      (@     `m@     @R@      @              :@     @R@      �?       @      G@      @     �m@      (@      f@      J@                       @      3@       @      �?      ;@      @      N@             �M@      5@      @      �?      4@     �M@      �?      @      I@      @     �S@      1@     �Q@     �A@              �?      (@      C@              @      ;@             �O@      "@     �I@      0@                       @      5@      �?       @      7@      @      .@       @      4@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJn*�ehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@%����@�	           ��@       	                    @�b�@S           ��@                           �?���ч%@�           <�@                          �1@b�HŖ@�            �v@������������������������       ���T�@:            �U@������������������������       �ؚߒbR@�            `q@                           �?�v~�	@�           �@������������������������       �ɋ�i��	@?           (�@������������������������       ���/~�@�            �k@
                          �4@��6��@�           ��@                          �1@o�n�@>           �@������������������������       �Lr��	 @�            �t@������������������������       �� B�@e           ��@                           @�`�`�@i            �e@������������������������       ��!�F��@1            �R@������������������������       �������@8            �X@                            �?/
�K�	@_           0�@                            �?��5�X	@E           ��@                           @V>�x�	@4           @}@������������������������       ���;	@           z@������������������������       ��=@�@            �I@                          �<@�!�`�@           �z@������������������������       �۾~,�{@�            0u@������������������������       ��mz��9@:            @U@                          �=@����@           ��@                          �7@}��tW@�           Ȇ@������������������������       ���>���@�            Pp@������������������������       ���EC\@*           @}@                           @�GEB�	@F            �]@������������������������       �&i��٘	@:            �X@������������������������       �l+�Y^�@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        >@     0r@     �@     �C@      L@     0|@     �T@     @�@      l@     ؈@      v@     �F@      *@     @\@      u@      2@      9@      j@      =@     ��@     �X@      @     �c@      1@      *@     �U@     �e@      .@      2@      a@      3@     �k@     �T@     �m@     �V@      $@              B@     �N@              �?      :@      @     �W@      3@     @Y@      5@      �?               @      6@                      @              <@      @      4@      @                      A@     �C@              �?      3@      @     �P@      ,@     @T@      2@      �?      *@     �I@      \@      .@      1@     �[@      .@     �_@     �O@     �`@     �Q@      "@      *@      F@      Q@      (@      (@      T@      $@     �Q@     �D@      Z@      K@      "@              @      F@      @      @      ?@      @     �L@      6@      ?@      0@                      :@     `d@      @      @      R@      $@     �{@      1@     @p@     @P@      @              7@      a@      @      @     �F@      @     Px@      ,@     @k@      L@      �?              @      E@              @      1@              e@       @     �T@      *@      �?              1@     �W@      @      @      <@      @     �k@      (@      a@     �E@                      @      ;@                      ;@      @     �I@      @      E@      "@      @              �?      4@                      "@      �?      7@      @      2@                               @      @                      2@      @      <@              8@      "@      @      1@     @f@     `n@      5@      ?@     @n@      K@      s@     @_@     �r@     �h@      <@      "@     �Y@     �\@       @      2@     �Z@      ?@     `b@     @T@     �b@      [@      1@      @      F@      N@      @      @      O@      6@      V@     �F@     �Q@     �F@      (@      @      B@     �L@      @      @     �M@      4@     @U@      >@      P@     �D@      @               @      @                      @       @      @      .@      @      @      @       @     �M@     �K@       @      &@     �F@      "@     �M@      B@     �S@     �O@      @      �?     �D@      G@       @      "@      F@      @      K@      :@     �Q@     �@@      @      �?      2@      "@               @      �?       @      @      $@      @      >@               @     �R@      `@      *@      *@     �`@      7@     �c@      F@     �b@      V@      &@      @     @P@      \@      @      @     �[@      3@     �b@      B@     �a@      Q@      &@              =@      I@       @      @      B@       @     �G@      @     �M@      7@      �?      @      B@      O@      @      �?     �R@      1@     @Y@      =@     @T@     �F@      $@       @      $@      0@      @      @      8@      @      &@       @      &@      4@               @      $@      0@      @      @      2@      @      @       @      @      1@                                       @              @              @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Ӿ3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��Z�X@�	           ��@       	                    @�r�/��@d           *�@                           �?���X��@�           �@                            �?~Y���@�            Pv@������������������������       ����5@J            @]@������������������������       �km� ��@�             n@                           @��h�2�@�           ��@������������������������       �ܪ��\�@�           X�@������������������������       ��@�f^�@             &@
                          �1@m΍��@�           h�@                           �?, h @�            Pw@������������������������       ����� @|            �h@������������������������       �ul��?p            �e@                           �?�'�-@�           (�@������������������������       �[��#T�?�             o@������������������������       �m6��}�@4           �~@                            �?�>}��@G           К@                            �?����@>           �@                           @��<~��@0           �~@������������������������       �-gm$F	@�             u@������������������������       ���j�>~@\             c@                          �<@���W@           @y@������������������������       �Ԭ�@Y�@�            �s@������������������������       ����*��@;            �U@                           �?q�NKf@	           ��@                           �?�O���@�            �i@������������������������       ���ĕz@;             V@������������������������       �C����@I            �]@                            @Ήx^�	@�           H�@������������������������       ��g�{�@z            `f@������������������������       �'��7Z	@           `{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �p@     �@      C@      N@     �{@     �U@     ��@     �i@     �@     Pw@      ?@      &@     @]@     �r@      .@      8@     �j@      A@      �@     �V@     �~@     �e@      .@      &@     @R@     `b@       @      3@     @b@      4@     �n@      R@     `m@     @X@      &@              8@      G@               @      ?@      �?     �Z@      (@      Y@      ?@      @              @      4@                       @              @@              G@      @                      4@      :@               @      7@      �?     �R@      (@      K@      8@      @      &@     �H@     @Y@       @      1@     �\@      3@      a@      N@     �`@     �P@       @       @     �H@     @Y@       @      1@     �\@      0@      a@     �M@     �`@     @P@      @      @                                      �?      @      �?      �?              �?      �?              F@     �c@      @      @     �P@      ,@      }@      2@     @p@      S@      @              @      G@               @      3@             @g@      @      V@      4@      �?              @      ;@               @      ,@             �Y@      �?      @@      1@                      @      3@                      @              U@      @      L@      @      �?             �B@     �[@      @      @     �G@      ,@     `q@      ,@     �e@      L@      @               @     �@@                      @      @      `@       @      N@      @                      =@     @S@      @      @      D@      $@     �b@      (@      \@      I@      @      &@     @c@     �m@      7@      B@     �l@     �J@     @s@     �\@     �t@      i@      0@      @     @S@     @^@      @      6@     �Y@     �@@      c@     @R@      f@     �\@      $@      @      C@      Q@      @      *@      O@      0@      X@     �C@     �U@     �K@      "@      @      @@     �E@              *@     �G@      "@      G@     �B@      N@     �B@      "@              @      9@      @              .@      @      I@       @      :@      2@               @     �C@     �J@       @      "@      D@      1@     �L@      A@     �V@      N@      �?      �?      =@     �F@       @       @      A@      *@     �H@      5@     �T@      @@      �?      �?      $@       @              �?      @      @       @      *@       @      <@              @     @S@     @]@      1@      ,@     �_@      4@     `c@     �D@     �c@     @U@      @              (@     �@@       @      �?      5@              L@      $@      K@      1@                      "@      2@       @      �?      (@              .@      @      ,@      &@                      @      .@                      "@             �D@      @      D@      @              @     @P@      U@      .@      *@     �Z@      4@     �X@      ?@      Z@      Q@      @       @      0@      2@      @      �?     �G@      @      <@      @      @@      1@      �?      @     �H@     �P@      &@      (@     �M@      ,@     �Q@      8@      R@     �I@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJcwn1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?De�m�N@�	           ��@       	                   �4@u-���@E           ��@                           @��X�,@           ��@                          �1@�9�F@�@�             u@������������������������       �Zy	���@E            �[@������������������������       ����x�	@�             l@                            �?&�WL(� @4           �~@������������������������       �Z�����?>             [@������������������������       �x�ӶAe@�             x@
                          @@@")�w��@D           p�@                            �?r�d�@1           H�@������������������������       ��:)h��@�            �k@������������������������       ���x�@�           P�@                           �?�8���l@            �B@������������������������       �bE��r @             2@������������������������       ��#p���@             3@                           �?9�i �{@s           >�@                          �<@��_�>x@q           ��@                          �2@��_u��@M            �@������������������������       �a����@x            @f@������������������������       �G��b�@�            �t@                            @���p`�@$             O@������������������������       �TfK@            �F@������������������������       ���ʙ��?             1@                          �:@�9};@           ��@                           @���W�@h           x�@������������������������       �r(�;��@'           ��@������������������������       ��qs{��@A           `�@                          �;@���2��	@�            0p@������������������������       �,M0MG@             F@������������������������       ����+��	@            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �p@     ��@      >@     �L@      ~@     �X@     H�@     @f@     ��@     �v@      >@       @     �Y@     p@      .@      ;@     �j@      E@      ~@     �N@     �s@      e@      &@      �?      >@     �\@      @      @     @Z@      $@     `s@      2@     �d@      Q@      �?      �?      7@     �O@      �?      �?     �O@      $@      Q@      *@      K@      C@      �?              @      ,@                      ,@      �?      C@      @      0@      1@              �?      0@     �H@      �?      �?     �H@      "@      >@      "@      C@      5@      �?              @     �I@       @      @      E@             @n@      @     �[@      >@                              @                       @             �M@              :@       @                      @      F@       @      @      A@             �f@      @      U@      6@              @     @R@     �a@      (@      7@     �[@      @@     �e@     �E@      c@     @Y@      $@      @      R@     �`@      (@      3@      [@      ;@     �e@     �E@      b@     �X@      $@       @      8@      ?@      �?              A@      @     �J@      "@      @@      ;@      @      �?      H@     @Y@      &@      3@     �R@      6@     �]@      A@      \@      R@      @      @      �?      &@              @       @      @                       @       @                              @              @      �?      �?                      @                      @      �?      @                      �?      @                       @       @              *@     `d@     u@      .@      >@     �p@     �L@     p~@     @]@     �@     �h@      3@             �E@     @W@      �?       @     �I@       @     `d@      0@     `d@     �B@      @             �A@     @U@      �?      �?      A@       @     �c@      (@     �c@      7@      @              (@      .@              �?      *@              T@       @      F@      &@                      7@     �Q@      �?              5@       @     �S@      $@     �\@      (@      @               @       @              �?      1@              @      @      @      ,@                      @       @              �?      "@              @      @      @      $@                      @                               @                      �?              @              *@      ^@     �n@      ,@      <@      k@     �K@     @t@     @Y@     pu@     �c@      0@      @      X@     �k@      *@      5@     �e@      D@     �r@     �R@      s@      \@      $@      @     �Q@     �b@      "@      5@     �a@      <@     �_@     @P@      b@     �S@      $@              :@     @Q@      @              A@      (@      f@      $@      d@     �@@              @      8@      8@      �?      @      E@      .@      5@      :@     �C@     �G@      @      �?      @                              @      �?      @      *@      @      @              @      5@      8@      �?      @      B@      ,@      ,@      *@     �@@      D@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @}����h@�	           ��@       	                    �?
S�p��@�           n�@                          �6@�-��F	@           ��@                           @P���E@<           ؋@������������������������       �7!x1��@�           �@������������������������       �pqHl�@�             k@                          �:@>^���	@�           p�@������������������������       ��8a�=	@           �z@������������������������       ���
�d�	@�            t@
                          �4@�~�ҩ�@�           p�@                           �?�?<��i@�             q@������������������������       �ڸ�%b�@<             W@������������������������       ������@z            �f@                            �?S;�@�            �s@������������������������       ����e:@w             e@������������������������       �E��J�@[            �b@                           �?;l�V&@5           H�@                           @�%���@5           P�@                           @�Qs��@|            �g@������������������������       �J{�"��@t             f@������������������������       ��0~�Ά@             *@                           @�;G�8D@�           h�@������������������������       �������@            {@������������������������       �������@�            `o@                            �?�9�/@            @�@                           @D"���}@{            �h@������������������������       �Pý��@S            �`@������������������������       �f���~@(            �O@                           �?�o�O_@�           �@������������������������       ��x��t@{            @g@������������������������       �X{��B@
           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     h�@     �A@     �J@     �}@      R@     H�@      m@     ؇@      v@     �A@      .@      l@     �t@      :@      F@     �u@     �J@     Pw@     `g@     �v@     �n@      =@      .@     @f@     �m@      9@     �C@     Pq@     �C@     @m@     `a@     �n@      g@      ;@      $@     @W@      `@      @      ,@     `a@      (@      f@     @Q@     �b@     �T@      "@      @      Q@     �W@      @      @     �W@      @     �b@     �C@     �`@     @P@      @      @      9@      A@               @     �F@      @      ;@      >@      1@      2@      @      @     @U@     �[@      2@      9@     @a@      ;@     �L@     �Q@     �W@     @Y@      2@              I@     �R@      $@      0@     @V@      &@      >@     �@@      L@     �F@      .@      @     �A@     �B@       @      "@     �H@      0@      ;@     �B@     �C@      L@      @              G@     @V@      �?      @     �P@      ,@     `a@      H@     �]@      N@       @              $@     �F@      �?       @      <@             �V@      .@     �N@      6@                      @       @                      &@              =@             �@@      @                      @     �B@      �?       @      1@             �N@      .@      <@      1@                      B@      F@              @     �C@      ,@     �H@     �@@      M@      C@       @              3@      5@              @      .@      (@      7@      1@     �D@      .@       @              1@      7@                      8@       @      :@      0@      1@      7@                     @W@     �l@      "@      "@     �`@      3@     ��@      G@     �x@     �[@      @              H@     �\@      @       @     �R@      @     Pu@      2@     �g@     �P@      @              0@      =@              �?      5@      @      N@      @     �@@      2@      �?              ,@      =@              �?      5@       @     �M@      @      @@      ,@      �?               @                                      @      �?      �?      �?      @                      @@     @U@      @      @     �J@      �?     �q@      ,@     �c@     �H@       @              2@     �G@              �?      ;@              h@       @     �Z@      @@       @              ,@      C@      @      @      :@      �?      V@      @      J@      1@                     �F@     �\@      @      �?      N@      (@     �q@      <@      j@     �E@      @              (@      8@      @              *@      @     @W@      @      >@      "@                      @      7@      �?              $@       @     �P@       @      3@      @                      @      �?      @              @      @      ;@      @      &@      @                     �@@     �V@       @      �?     �G@      @     @h@      6@     @f@      A@      @              @     �B@              �?      @      @     @R@      @     �G@      @      �?              ;@      K@       @              D@      �?     @^@      .@     ``@      ?@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�ӱ�5@�	           ��@       	                    �?��z8/@           x�@                           �?m��F8@3           �~@                          �4@��@�             m@������������������������       �d�����@A             X@������������������������       �I���M@U             a@                            @<Z���@�            pp@������������������������       �vx����@e            `c@������������������������       �B��?�@8             [@
                            @�<�1�@�           x�@                          �8@ŏ�0�C@y           ��@������������������������       �i�3|@@           �@������������������������       ���p�@9            �U@                          �7@M:r1��?X            @c@������������������������       �v.ꪈ�?=            �Z@������������������������       ����?             H@                           @�Fi�3@�           ֤@                           @8~��~	@�           4�@                          �3@����	@u           `�@������������������������       ���Q�@�            �q@������������������������       �}����7	@�           ��@                           �?<%C�3�	@t           �@������������������������       �Yb-�� 
@            {@������������������������       �����+@[            �a@                           !@���@�           x�@                           @�Jߙ��@�           @�@������������������������       �M�c׉�@�           ؈@������������������������       �ԩ<�@�            Ps@������������������������       �JE}�u) @             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@      r@     ��@      =@     �J@     @}@     �U@     ��@     �j@     h�@     pt@      @@             �V@     @f@      �?      "@     �X@      (@     �|@     �B@     �r@     �N@      @             �I@     @V@               @     �N@      @      [@      5@     �\@      B@      @              4@     �E@              @      A@      @      G@      0@     �G@      0@                      @      6@                      (@      @      :@      @      3@      @                      1@      5@              @      6@              4@      (@      <@      "@                      ?@      G@              �?      ;@              O@      @      Q@      4@      @              0@      5@              �?      .@              A@      @     �J@      "@      @              .@      9@                      (@              <@       @      .@      &@                     �C@     @V@      �?      �?      C@      "@     �u@      0@     �f@      9@       @              >@      U@      �?              A@      "@     �p@      &@      a@      8@       @              >@      Q@      �?              ?@      @     �m@      @     @]@      1@       @                      0@                      @      @      =@      @      3@      @                      "@      @              �?      @             �T@      @      G@      �?                      @      @              �?                      M@              A@      �?                       @                              @              9@      @      (@                      2@      i@     �v@      <@      F@     w@     �R@     @�@     @f@      �@     �p@      ;@      1@     @a@     �j@      8@     �A@     p@      L@      j@     �b@     �o@     `e@      9@       @      T@     @_@      0@      3@      e@      B@     �`@     �Q@      g@      ^@      (@      @      0@     �E@       @      @      =@      @      O@      4@     �L@     �D@              @      P@     �T@      ,@      *@     `a@      ?@      R@      I@     �_@     �S@      (@      "@      M@     @V@       @      0@     @V@      4@     �R@     @T@     @Q@     �I@      *@      "@     �G@     �Q@      @      (@      S@      1@      H@     �J@      C@      F@      *@              &@      3@      �?      @      *@      @      :@      <@      ?@      @              �?      O@     �b@      @      "@      \@      3@     �u@      ;@     pr@     �W@       @      �?     �M@     `b@      @      "@     @[@      *@     �u@      ;@     `r@     �W@       @      �?     �A@     �Z@      �?      @     �Q@      @     0q@      .@     �k@     �N@       @              8@     �D@      @      @     �C@       @     @Q@      (@     @R@      A@                      @      �?                      @      @                      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�BhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�s7?�)@�	           ��@       	                    �?��ռRJ	@           D�@                           �?s�L<u@%           �|@                            @��]�@@s            `g@������������������������       �x��"B@T            �a@������������������������       �B����=@            �G@                          �5@�:�@�             q@������������������������       �2Hii;@T             `@������������������������       �z-�p�@^            @b@
                           �?e,�
�	@�           �@                           �?�<޹2#@;            @X@������������������������       ���^�q�@             9@������������������������       �i^�P0�@.             R@                          �:@�1��	@�           ��@������������������������       ���~�(t	@           ��@������������������������       ���۩��	@�             n@                           �?����e�@�           �@                           @�_]���@�           p�@                           �?�)K&s@r            �f@������������������������       � @�?��@>            @X@������������������������       �3�<�j�@4            @U@                            �?N� � @e           ��@������������������������       �~*y�L�?K            �^@������������������������       �,�2��Q@           �{@                          �3@n8xٽ@�           (�@                           @_�e�?@}           ��@������������������������       ���UM@;             W@������������������������       ������B@B           ��@                           �?��Am�@V           ��@������������������������       �,.�0�@$             L@������������������������       ��a<ɖ�@2           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `p@     p�@     �B@      K@      }@      S@     D�@     �h@     ��@     �w@      ?@      2@     @b@     `k@      7@     �B@     @o@     �H@     �m@     @`@     �p@     �j@      7@      @      D@      P@      @      @      Q@      @     @X@      ;@      U@     �O@      @      @      0@      1@                      8@             �I@      @      I@      5@      �?      @      *@       @                      7@              ?@      @     �C@      3@      �?              @      "@                      �?              4@      �?      &@       @                      8@     �G@      @      @      F@      @      G@      7@      A@      E@       @              4@      &@       @       @      1@       @     �B@      @      .@      ,@      �?              @      B@      �?      @      ;@      �?      "@      0@      3@      <@      �?      .@     �Z@     `c@      4@      ?@     �f@      G@     �a@     �Y@      g@     �b@      4@      @      @      "@              @      4@      @              (@      8@      .@      �?       @      �?      @                      @      @               @              @              �?      @      @              @      .@      @              $@      8@       @      �?      (@     �Y@     @b@      4@      <@     @d@      D@     �a@     �V@      d@      a@      3@      @     �S@      ^@      .@      7@      `@      ;@      _@     @Q@     �_@     �U@      1@      "@      8@      :@      @      @     �@@      *@      2@      6@     �A@     �H@       @       @      ]@     0s@      ,@      1@      k@      ;@     �@     @Q@     H�@     �d@       @              A@      Y@      �?       @      G@      @     @u@      $@     �f@      =@      @              &@      0@              �?      6@      �?      R@      @     �F@      @      @              @      &@              �?      0@      �?     �B@      @      2@      @                      @      @                      @             �A@      �?      ;@      @      @              7@      U@      �?      �?      8@       @     �p@      @      a@      6@      �?                      ,@      �?              "@      �?     �R@      �?      4@       @                      7@     �Q@              �?      .@      �?     @h@      @      ]@      4@      �?       @     �T@     �i@      *@      .@     @e@      8@     �|@     �M@     @w@      a@      @              8@     @X@      �?      @      E@      �?     @n@      1@     @c@     �F@                      @      0@               @      "@      �?      A@      @       @      "@                      2@     @T@      �?       @     �@@              j@      $@     @b@      B@               @      M@     �[@      (@      &@      `@      7@     �k@      E@     @k@     �V@      @       @      @       @              @      @      @      �?      @      2@      @                     �J@     �Y@      (@      @      _@      3@     `k@     �C@      i@     @U@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ`�u}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @���[w%@�	           ��@       	                    �?><E�@�           h�@                           �?'D�"
@�           X�@                           �?��Ae�@7           �}@������������������������       �y�Hm$<@�            �k@������������������������       ��s�T�R@�            �o@                            �?�8�V@v            �i@������������������������       ���ؒ���?&            @R@������������������������       ��$�g�@P            �`@
                           �?�ZRmX	@�           $�@                           �?��L(��	@�           �@������������������������       ���aE@            z@������������������������       �x��B�	@�            �@                           �?����I@           0|@������������������������       ���ZI!@e             e@������������������������       �N{s��@�            �q@                            �?S�C�@'           T�@                           @~Erz2C@S           ȍ@                          �7@)�I�
@H           @�@������������������������       �H�I�@�           x�@������������������������       ���(�9@x             g@������������������������       ��65�@             1@                          �4@�;.=@�           ��@                          �1@�|a�w @�            �x@������������������������       ��q�]�_�?X            �a@������������������������       �x���@�            �o@                          �9@$�s��^@�            @u@������������������������       ����O�@�            �m@������������������������       ��yHh�"@C            @Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     �r@     `�@      =@     �K@     0z@     �R@     ��@      l@     �@     x@      =@      ,@      k@     0s@      7@      D@      r@      K@     Py@      g@     �y@      p@      <@      �?     �R@     �T@       @      @     �O@       @      h@     �B@      c@      P@      @      �?     �M@     �P@       @      @     �H@       @      [@      =@     @X@     �I@      @      �?      ;@      =@       @      @      :@       @     �G@      5@     �A@      9@      �?              @@      C@                      7@             �N@       @      O@      :@      @              .@      0@                      ,@             @U@       @      L@      *@                              @                      @              C@              9@       @                      .@      &@                      &@             �G@       @      ?@      &@              *@     �a@      l@      5@     �@@     `l@      J@     �j@     �b@      p@      h@      8@      *@     �Z@     �b@      ,@      7@     �d@      D@     ``@     @[@     �e@     @b@      6@      @      5@      P@      @      @      O@      "@     @S@     �C@     �P@     �N@      @      $@     @U@      U@      &@      0@     @Z@      ?@      K@     �Q@      [@     @U@      1@             �B@      S@      @      $@      N@      (@     @T@     �C@     @T@      G@       @              ,@      =@      @      �?      7@      @      6@      ,@      B@      5@       @              7@     �G@      @      "@     �B@      "@     �M@      9@     �F@      9@               @     �S@      k@      @      .@      `@      5@     p�@      D@     �x@      `@      �?             �J@     @`@      @      @     �Q@      .@     Pu@      6@      l@      V@                     �G@     @`@      @      @     �Q@      (@     @u@      5@     �k@      V@                      ?@     �Z@      @      @     �J@      @     0s@      ,@     �e@      J@                      0@      7@              �?      1@      @     �@@      @      G@      B@                      @                      �?              @      �?      �?      @                       @      :@     �U@       @      $@     �M@      @     �s@      2@     �d@     �D@      �?              (@      G@              @      4@      @     @j@       @     �S@      "@                      @      *@                      &@             �R@      �?      C@                              "@     �@@              @      "@      @      a@      @     �D@      "@               @      ,@     �D@       @      @     �C@       @     �Y@      $@      V@      @@      �?       @      $@      ?@      �?              >@       @      S@       @      L@      <@      �?              @      $@      �?      @      "@              ;@       @      @@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�F�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?	D�ЈY@�	           ��@       	                    �?��0/՟@4           �@                           �?>=�z�L@<           }@                            @�{h�ԧ@z            `e@������������������������       �ǵ�e0@Z            @`@������������������������       ��c��@             �D@                            @t�ML�@�            `r@������������������������       ���)F@j            �c@������������������������       �X5�l�|@X             a@
                           �??���@�           H�@                           @(�B�b�@            �|@������������������������       ��.i�g�@s            �g@������������������������       � ��:tG�?�            �p@                          �8@h?�@�            �u@������������������������       �O���� @�            q@������������������������       �N�Zyo@-             S@                           @�_�*bD@�           ��@                          �1@d�Gt @�           �@                           @�,[S��@�            v@������������������������       �1Fgj�@              L@������������������������       ��X���M@�            �r@                          �9@?�`��z@�           ��@������������������������       ��J��@�           ��@������������������������       �a�[�\	@           �z@                           @G�Sk	@�            Pt@                           �?�_8y�[
@�            �i@������������������������       ��'���	@.            @Q@������������������������       ��A�U�	@R            �`@                          �:@(FZ�7@D            @^@������������������������       �m�R���@9            �X@������������������������       �>Gzuw�?             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      r@     ��@      ?@      K@     �{@     �S@     p�@     �k@     Ј@     �w@     �B@       @     �U@     �h@       @      "@     �Z@      0@     �|@      C@     @q@     @S@      @       @     �L@     �U@      �?      @     �G@      @      W@      ;@      W@      G@      @       @      5@      6@                      5@             �F@      @     �B@      1@      �?       @      2@      ,@                      3@              ;@      @      =@      0@      �?              @       @                       @              2@      �?       @      �?                      B@      P@      �?      @      :@      @     �G@      6@     �K@      =@      @              6@      <@      �?      @      $@       @      5@      (@     �A@      2@      @              ,@      B@               @      0@       @      :@      $@      4@      &@                      =@     �[@      �?      @      N@      (@     �v@      &@      g@      ?@      �?              0@     �P@              @     �D@       @     �l@      @     �R@      2@                      &@      >@               @      8@       @     �Q@      @      >@      &@                      @     �B@              �?      1@             �c@      �?      F@      @                      *@     �E@      �?              3@      @     `a@      @     �[@      *@      �?              *@     �A@      �?              *@             �]@      @     �T@      @                               @                      @      @      4@       @      <@      @      �?      .@     �i@     �v@      =@     �F@     @u@     �O@     �@     �f@     0�@     �r@      ?@      "@     `f@     ps@      9@     �E@     �r@     �J@     @      c@     p}@     p@      3@              (@      L@               @      6@             �]@      3@      W@      @@                      @      @                      �?              8@       @      "@      @                      @     �J@               @      5@             �W@      &@     �T@      :@              "@     �d@     �o@      9@     �D@     @q@     �J@     �w@     �`@     �w@      l@      3@      @     �]@      k@      3@      A@      k@     �A@      t@     @T@     t@     `c@      ,@      @     �H@     �C@      @      @     �M@      2@     �M@      J@      M@     �Q@      @      @      9@     �K@      @       @      E@      $@      I@      >@     �G@      E@      (@      @      3@      A@      @       @      ;@      $@      8@      8@      0@      ;@      (@              "@      @       @      �?      &@      @      @      $@      @      (@      @      @      $@      <@      �?      �?      0@      @      5@      ,@      &@      .@      @              @      5@      �?              .@              :@      @      ?@      .@                       @      1@      �?              @              :@      @      <@      ,@                      @      @                      &@                              @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��vyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �7@1$�:�s@�	           ��@       	                   �1@[�>@�           ��@                           @����5�@�           ��@                           @��|<�@�            �r@������������������������       ��qˌm�@�            @q@������������������������       ��
E�� @	             4@                           @�s[#Rt @�            �t@������������������������       ��JY�Ƿ�?l            �d@������������������������       �����r� @s             e@
                          �4@� yq�@#           ��@                            @%��T@�           @�@������������������������       ��B���@"           �@������������������������       ����?@�            �t@                           @���[b@6           ��@������������������������       ��te�	�@[           Ȁ@������������������������       �7EY�@�            Pv@                          �;@ʃ�eP	@�           �@                           @dd�X@�@�           @�@                            �?���=�K@�           p�@������������������������       ��^���]	@q            `f@������������������������       ��Pϟ�l@%           �{@                            �?�s^��|@:            �V@������������������������       ���9=^W@"            �I@������������������������       ���6�κ@            �C@                          �?@;7o��	@           �{@                          �>@����f	@�            pu@������������������������       ���M=	@�            �q@������������������������       ��M���@#             O@                            �?3n�@A             Z@������������������������       �	��N�@             ?@������������������������       �L���@/            @R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     Pq@     0�@      ?@     �J@     �@     @V@     �@     �j@     P�@     �v@      B@      (@     �e@     �x@      0@      8@     Pt@     �I@     0�@      _@     ��@     �j@      ,@              7@     �U@      �?      @     �P@      @      p@      9@     �^@     �D@                      *@     �K@      �?      �?      G@      @      V@      6@      E@      9@                      (@     �K@      �?      �?     �C@              V@      6@     �B@      5@                      �?                              @      @                      @      @                      $@      ?@              @      4@              e@      @      T@      0@                      "@      &@                      (@              Y@      �?      7@       @                      �?      4@              @       @              Q@       @     �L@       @              (@      c@     �s@      .@      3@     0p@      H@     0�@     �X@     �{@     �e@      ,@      @     @T@     `e@      @       @     �`@      2@     @v@      P@      q@     �Y@      $@             �L@     @`@      @      @     �V@      &@     @q@     �I@     �g@     @S@      @      @      8@     �D@       @      @      F@      @      T@      *@      U@      :@      @      @     �Q@     �a@      "@      &@      _@      >@     @l@     �A@     �d@     �Q@      @      @     �O@      W@      @      $@      U@      5@     �T@     �@@     @W@     �F@      @               @      I@      @      �?      D@      "@     �a@       @     @R@      9@      �?      &@     �Y@     �b@      .@      =@     �f@      C@     �c@     @V@      k@     �b@      6@      �?     �H@     �W@      @      0@      ]@      7@      \@     �O@      c@      P@      .@              C@     @T@      @      0@     �Z@      3@     �X@      I@     �`@      O@      &@              1@      1@              "@      3@      "@      :@      2@      B@      5@      @              5@      P@      @      @      V@      $@      R@      @@     �X@     �D@      @      �?      &@      ,@      �?              "@      @      ,@      *@      1@       @      @              @      @      �?              @       @      @      "@      0@       @              �?      @      "@                      @       @      "@      @      �?              @      $@     �J@      L@      "@      *@     @P@      .@      F@      :@      P@     @U@      @      @      9@     �I@      @      $@     �J@      ,@      C@      1@      I@     �P@      @      @      9@      G@      @      @      D@      *@      >@      *@     �E@     �I@                              @              @      *@      �?       @      @      @      0@      @      @      <@      @       @      @      (@      �?      @      "@      ,@      2@       @              @      �?                       @              @      @       @      @       @      @      7@      @       @      @      $@      �?      �?       @      (@      &@        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�\_\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?U~Ù,L@�	           ��@       	                   �3@�>��V.@+           d�@                            �?��s��@�           Ȅ@                           @��h�@d            `d@������������������������       ��Y�Tَ@<            �X@������������������������       ���;��S�?(            @P@                          �1@��@2R@;           `@������������������������       �l�I�B�@�            �l@������������������������       �� :��@�            �p@
                           �?C�ķ#�@�            �@                           �?��
��D@�            �v@������������������������       �Y��4Z�@^            �c@������������������������       �pı_�@�            �i@                           @��	@�           ��@������������������������       ���K_.	@h           ��@������������������������       �����@;             Y@                           @���M@|           `�@                           �?�o�W�@a           ��@                          �<@�M��ٰ@�            �v@������������������������       �l��O'�@�            t@������������������������       ���SA��@             F@                           �?��i3�\	@~           �@������������������������       ��'n�	@�           �@������������������������       ������@�            �q@                          �7@��CL�@           �@                            �?=󚊍\@�           ��@������������������������       ��rW�@�            `u@������������������������       �a]�VMI@�            �q@                            @|����@�            �i@������������������������       �LW5x��@j            �c@������������������������       ��.u��@             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     @q@     �@     �B@      O@     {@     �W@     4�@     �i@     ��@     pu@      9@      *@     �]@      l@      1@      ?@     �f@      F@     �@      S@     �s@     `b@      (@      @      3@      R@       @      @     �Q@      @     �q@      5@     �`@     �H@       @              �?      7@              �?      5@       @     �P@      &@      9@      $@       @              �?      1@                      *@       @      >@      &@      ,@       @       @                      @              �?       @             �B@              &@       @              @      2@     �H@       @      @     �H@      @     �j@      $@     @[@     �C@               @       @      8@       @      @      6@             �\@      �?      D@      ,@              @      $@      9@                      ;@      @      Y@      "@     @Q@      9@               @      Y@      c@      .@      ;@     �[@     �C@     �l@     �K@     �f@     �X@      $@      �?      >@     �K@       @      (@      @@      @      ^@      ,@     �P@      7@       @      �?      3@      =@       @      &@      ,@       @      6@      &@      A@      "@       @              &@      :@              �?      2@      @     �X@      @     �@@      ,@              @     �Q@     �X@      *@      .@     �S@      A@      [@     �D@     @\@     �R@       @      @     �L@     �U@      *@      .@      N@      =@     �W@      9@     �Y@     �Q@      @      �?      *@      &@                      3@      @      ,@      0@      &@      @      @      *@     �c@     t@      4@      ?@     �o@      I@     x�@      `@      �@     �h@      *@      *@     �]@     �i@      2@      >@     @h@     �A@     �l@     @Z@     Pr@      a@      (@              >@      M@               @     �B@              X@      $@     �Y@      :@      @              9@     �I@                      >@             @W@      @      X@      2@       @              @      @               @      @              @      @      @       @      �?      *@      V@     �b@      2@      <@     �c@     �A@     �`@     �W@     �g@     �[@      "@      *@      R@      V@      .@      3@      [@      ;@     �R@      R@     `c@     �U@      "@              0@     �N@      @      "@     �H@       @     �M@      7@     �A@      8@                     �C@     �\@       @      �?      M@      .@     �r@      7@     �k@     �M@      �?              ;@      X@      �?      �?      4@      "@     �n@      &@     @f@      C@      �?              3@     �I@      �?      �?      ,@      �?     �^@      @     @X@      @@                       @     �F@                      @       @     @^@       @     @T@      @      �?              (@      2@      �?              C@      @      K@      (@     �F@      5@                       @      2@                      9@      @     �D@      "@     �A@      1@                      @              �?              *@              *@      @      $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ophG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @N���e@�	           ��@       	                   �4@��� �@�           ֥@                           @6��n/�@=           ��@                           �? %/p�U@_           ��@������������������������       ���J���@w            @g@������������������������       �!��[�,@�            pw@                          �1@��k��@�           ��@������������������������       �inb�0��?�            �p@������������������������       ��9�)7d@%           �~@
                          �<@怓�F@�           �@                            �? ({z��@           ��@������������������������       ���}�k�@8           �@������������������������       ���a�&@�           h�@                           �?ގs���@�            �j@������������������������       �Я�h��@-            �S@������������������������       ��\"�@]             a@                           @��6L@�           x�@                          �1@�����)	@            �@                          �0@JlɄ	@>             X@������������������������       ���&x�@             8@������������������������       �v�T_��@0             R@                           �?��U-:	@�            �@������������������������       �V�n���@s             h@������������������������       �EC��a�	@b           �@                           @{d`C�l@�            �q@                           @������?h             d@������������������������       �9��<��?/            �R@������������������������       �lx 8��?9            �U@                           @��dOl�@R            �^@������������������������       ����W�7�?'            �M@������������������������       �X�Ч�>@+            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �r@     ��@     �@@      L@     �}@     @S@     ��@     �l@      �@      u@      :@      $@     �h@     �x@      1@     �A@     @t@     �N@     p�@     @d@     ��@     �m@      0@             �P@     �e@      "@      $@     �_@      ,@      ~@     �N@      q@     @X@      @             �F@     @P@      @      @     �U@      (@     `b@      F@      W@     �K@      @              &@      5@              �?      9@             �P@      $@     �B@      *@       @              A@      F@      @      @     �N@      (@     @T@      A@     �K@      E@      @              5@      [@      @      @     �D@       @     �t@      1@     �f@      E@                      �?      :@               @      (@             �b@      @     �M@      ,@                      4@     �T@      @      @      =@       @      g@      *@     �^@      <@              $@     �`@     �k@       @      9@     �h@     �G@     �p@     @Y@     �s@     `a@      "@      $@     �Z@     @h@      @      6@     �d@     �D@     �o@     �S@     �q@     �W@      @      @     �L@     �P@      @      *@      P@      .@     @Y@     �A@     @Y@      F@      @      @      I@     �_@      @      "@      Y@      :@     @c@     �E@     `f@     �I@       @              9@      ;@      �?      @     �@@      @      *@      7@      C@      F@       @              ,@      1@                      @      �?      @      "@      $@      0@                      &@      $@      �?      @      :@      @      "@      ,@      <@      <@       @      0@     �Y@      e@      0@      5@      c@      0@     �m@     �P@      j@     �Y@      $@      0@     @W@     @b@      .@      2@      `@      ,@      ^@      P@     ``@     @T@      $@              @      "@       @       @      "@              @@      .@      4@       @                              �?               @      @              @      @      @                              @       @       @              @              =@       @      ,@       @              0@      V@      a@      *@      0@     �]@      ,@      V@     �H@     �[@     �S@      $@              3@      G@       @      �?      9@              @@       @     �C@      5@              0@     @Q@     �V@      &@      .@     �W@      ,@      L@     �D@      R@      M@      $@              $@      6@      �?      @      9@       @     �]@      @     @S@      5@                      @      "@                      &@      �?     �P@       @      N@      @                      @      @                              �?     �@@       @      <@                               @      @                      &@              A@              @@      @                      @      *@      �?      @      ,@      �?     �I@      �?      1@      1@                      �?      �?                      @             �C@      �?       @      @                      @      (@      �?      @       @      �?      (@              "@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ|�ZUhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�6!�a@�	           ��@       	                   �<@^ti� r@           �@                           �?s�赛@�           ��@                          �0@q=��@           �z@������������������������       ��!�:f��?             5@������������������������       �`A����@           Py@                            �?�[��H@�           ؅@������������������������       �������?z            �f@������������������������       ��i��M@S            �@
                          �>@d3���@=            @X@                            �?)P�$X@"            �K@������������������������       ��[���@             (@������������������������       ��Q��@            �E@                           @uH�Y�2@             E@������������������������       �^~m��D@             ?@������������������������       �lofON@             &@                          �5@#��t�Q@�           �@                           @�qv2O�@m           ؕ@                          �2@Z�	}�@�           @�@������������������������       ���c��@�            �s@������������������������       ��{�n[@           �z@                           �?��o�g�@�           p�@������������������������       ��Է+@�            �t@������������������������       ���Qj�@�            @t@                           @�ICA@s	@'           4�@                          �;@� [V0�	@           �@������������������������       �1@|��y	@q           ��@������������������������       �bt��
@�             n@                          �6@
�}�	@!           �|@������������������������       ���r�S�@5            @U@������������������������       ��V��(�@�            Pw@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �t@     `�@      ;@      K@     �}@      R@     p�@     �l@     Ȉ@     �u@      B@      �?     �S@     @d@      @      @     �\@      "@     �z@      F@     �r@     @R@      @      �?     �P@     �b@      @      @     �X@       @     @z@      ?@      r@      K@      @      �?      D@     �P@               @      P@       @     �W@      4@     �Y@      >@       @              �?                              &@              @               @      �?              �?     �C@     �P@               @     �J@       @     @V@      4@     @Y@      =@       @              ;@     @T@      @      �?     �A@      @     Pt@      &@      g@      8@      �?              �?      4@      @      �?      @      @      Y@              C@      "@                      :@     �N@                      <@       @      l@      &@     `b@      .@      �?              (@      ,@              @      .@      �?      @      *@      &@      3@       @              @       @              �?      @              @       @       @      1@       @                      @                      @                               @      �?       @              @      @              �?       @              @       @      @      0@                      @      @               @      $@      �?              &@      @       @                      @      @               @      @                       @       @                                      �?                      @      �?              @      �?       @              ,@     �o@     �x@      8@      H@     �v@     �O@     �@     `g@     �~@     @q@      ?@      @     @U@     `j@      "@      2@     `e@      8@     0w@     @T@     s@      ]@      @      @      L@      \@      @      .@      ]@      3@     �a@      R@     �`@      Q@       @      �?      7@     �G@      �?      @     �@@       @     �S@      B@      L@      ?@      �?       @     �@@     @P@      @      (@     �T@      1@     �O@      B@     �S@     �B@      �?              =@     �X@      @      @     �K@      @     �l@      "@     @e@      H@       @              3@     �I@      @       @      C@       @      Z@       @     �R@      :@      �?              $@      H@              �?      1@      @     @_@      �?      X@      6@      �?      &@      e@     �f@      .@      >@     �g@     �C@      f@     �Z@     �g@      d@      ;@      $@     @]@     �]@      "@      5@     �_@      A@      R@     �U@     �V@     @^@      ;@       @      V@     �U@      @      .@      Y@      9@     �K@     �P@     �O@     �Q@      5@       @      =@     �@@      @      @      ;@      "@      1@      4@      <@     �I@      @      �?     �I@      P@      @      "@      O@      @      Z@      3@     �X@     �C@                      $@      @      @              .@              @@              (@      @              �?     �D@     �M@              "@     �G@      @      R@      3@     �U@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ5�N-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?<�3���@�	           ��@       	                    �?�����@�           ��@                          �<@��1�d3@�           ��@                           �?TW�C�@s           ��@������������������������       ��*z���@{             i@������������������������       �Z~2��7@�            �x@                           �?��K�=2@             F@������������������������       �@�lB��?            �@@������������������������       �@	B0f@
             &@
                          �6@��<@`           ��@                           �?ʼ����@�            �w@������������������������       �A�y�q@M            �]@������������������������       ��C��dt @�             p@                           �?$<G��@v            @g@������������������������       �����8�@B            �\@������������������������       �^ �3a�@4            �Q@                           @�a�1�n@�           2�@                           �?���e$B	@�           ��@                           �?�5(e��	@�           Б@������������������������       ��tA*�@           �{@������������������������       �j[NW��	@�           ��@                           �?[�tջu@           �|@������������������������       �jZp
�@             D@������������������������       �;�v�
@           0z@                           @K��0-@�           h�@                          �1@N��(E@�            �@������������������������       ���[*b2�?]            `b@������������������������       ��>h��G@�           h�@                           @��q��f@�            �s@������������������������       �e�b�@�            0q@������������������������       ���Nb	@            �C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     (�@      ?@     �O@     |@     �U@     X�@      l@     @�@     `x@     �@@             �T@     @e@       @      @     �V@      $@      z@      @@     0q@     �W@      (@              C@     �X@      @      @      G@       @     �o@      (@     @_@      G@       @             �B@     @V@      @       @      F@      @     �n@      &@     �]@      =@       @              3@     �@@      @              6@       @      K@      "@     �C@      *@       @              2@      L@               @      6@      @      h@       @      T@      0@                      �?      "@               @       @      �?      @      �?      @      1@                              "@               @       @               @               @      0@                      �?                                      �?      @      �?      @      �?                      F@      R@      �?      @     �F@       @     �d@      4@     �b@     �H@      $@              :@      F@               @      1@             @a@      &@     �\@      6@       @              (@      5@               @      *@              7@      @      ?@      *@                      ,@      7@                      @             �\@       @     �T@      "@       @              2@      <@      �?      �?      <@       @      <@      "@      B@      ;@       @              0@      2@              �?      3@              ,@      @      .@      2@      @               @      $@      �?              "@       @      ,@       @      5@      "@      �?      5@     �m@     �w@      7@      L@     `v@     @S@     H�@      h@     P@     pr@      5@      3@     `d@     �m@      (@     �C@     �n@      M@      l@     @c@      m@     �h@      .@      3@     ``@     �b@      (@      >@      g@      F@     �`@     �\@     �c@     �b@      ,@      @      ;@     �Q@      �?      .@     �Q@      *@     @Q@     �F@      O@     �N@      @      0@      Z@     �S@      &@      .@     �\@      ?@     @P@     �Q@     �W@     @V@      &@              @@     @V@              "@     �N@      ,@     �V@     �C@     �R@     �H@      �?              @      @              @      $@      �?       @      @      @      @                      <@     @U@              @     �I@      *@      V@      A@     �Q@      F@      �?       @     @R@     �a@      &@      1@      \@      3@     �t@     �C@     �p@      X@      @       @     �L@     @Z@      �?      "@     �T@      &@     pp@      6@     �g@     �J@      @              @      .@                      @             @R@              H@      @               @      K@     �V@      �?      "@     �S@      &@     �g@      6@     �a@     �H@      @              0@      B@      $@       @      >@       @     �P@      1@      T@     �E@                      ,@      @@      @      @      9@      @     �N@      (@     �R@     �C@                       @      @      @      �?      @      �?      @      @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJZdhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����c@�	           ��@       	                    �?(`�Q	@           H�@                           �?_'oS�@.           }@                            �?��9�h@�             k@������������������������       �:4W�FX@C             [@������������������������       ��}ۣk@L            @[@                          �5@*X�І@�             o@������������������������       �n��ݢ�@T            @a@������������������������       ���oϦw@K            �[@
                           �?(��I(�	@�           �@                          �1@��.���@           {@������������������������       �|�[90@!             O@������������������������       ��%�'[�@�            0w@                          �6@
���hH
@�           ��@������������������������       ����o�@�            v@������������������������       ���CW��
@�            �v@                           �?��9��@�           �@                          �;@�ٚ�tD@�           8�@                            �?�1���@�           ��@������������������������       �n�F�1@�            pw@������������������������       �YC{V֥ @�            pt@                           @����S�@            �D@������������������������       �b�H�@             4@������������������������       ��� ���?             5@                           �?��z�@�           @�@                            @��6���@G             \@������������������������       ���S�b@9            �U@������������������������       ���a��#@             :@                          �4@9����@�           ��@������������������������       �埽÷@�           X�@������������������������       ��w���@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     @�@      =@     �J@     �|@     @S@     ��@      p@     p�@     pu@      A@      3@     @e@      m@      2@     �A@     @p@      F@      n@      c@     �n@     �e@      <@             �I@     @S@       @      @     �L@      @      [@      >@     @W@     �B@       @              9@      >@       @      @      >@      @     �I@      1@      A@      5@                      .@      3@              �?      2@              7@      $@      $@      (@                      $@      &@       @      @      (@      @      <@      @      8@      "@                      :@     �G@              �?      ;@             �L@      *@     �M@      0@       @              (@      <@              �?      "@              F@      @      A@      @                      ,@      3@                      2@              *@      $@      9@      "@       @      3@     �]@     `c@      0@      >@     `i@     �D@     �`@     �^@      c@      a@      :@      @      <@     �N@      �?      (@     @S@      "@     �O@      M@      O@      J@      @              @      @                      @       @      :@              $@       @              @      6@     �L@      �?      (@     �Q@      @     �B@      M@      J@      F@      @      .@     �V@     �W@      .@      2@     �_@      @@     @Q@      P@     �V@     @U@      4@      @      I@     �F@      @      @     �O@      @      D@      <@     �N@      D@      @       @     �D@     �H@      (@      .@     �O@      :@      =@      B@      >@     �F@      *@      �?     �_@      t@      &@      2@     �h@     �@@      �@      Z@     ��@      e@      @             �A@     �U@              @     �E@       @     0u@      1@     �e@     �A@      �?              ;@      U@              @     �C@      @     0t@      (@     �e@     �@@                      ,@     �N@              @      <@       @     @c@       @     �V@      3@                      *@      7@               @      &@      @      e@      $@     @T@      ,@                       @       @                      @       @      0@      @      �?       @      �?               @      �?                       @               @      @              �?      �?                      �?                       @       @      ,@              �?      �?              �?      W@     @m@      &@      (@     `c@      9@     {@     �U@     �v@     �`@      @      �?      @      1@              @      0@       @      (@      1@      5@      1@              �?      @      *@               @      ,@      �?      $@      "@      4@      &@                              @               @       @      �?       @       @      �?      @                     �U@      k@      &@       @     `a@      7@     Pz@     �Q@     `u@     @]@      @              >@      ^@      "@      @      J@       @     @o@      =@     �e@      E@                     �L@     @X@       @       @     �U@      5@     `e@     �D@     �d@     �R@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��dshG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?a�@�	           ��@       	                    @i����@�           ��@                          �;@;�K�@�           ��@                          �7@�+9�@Z           X�@������������������������       ����S	o@           y@������������������������       ������@L            �^@                           �?���H0@7            @T@������������������������       �7Q/���@+             P@������������������������       ��o���@             1@
                          �4@=	CE~@e           h�@                           �?����?�            `v@������������������������       �d�ɛr�?�            �j@������������������������       �;�ǤL�?W             b@                            @QR���[@�            �l@������������������������       �����@r            `f@������������������������       ���* W�?             J@                            @g���f@�           @�@                          �4@+��@�           ��@                          �1@������@           ��@������������������������       ��w-RUW@�            �o@������������������������       �.P����@u           ؂@                          �8@��	&A	@�           4�@������������������������       ���o8��@}           `�@������������������������       �W��e�_	@/           ~@                           @�D�9��@�           ؇@                          �9@���Ѥz	@�           P�@������������������������       ��wDQ�@&           0|@������������������������       ���o��	@_            �d@                           @ ��@d             b@������������������������       �f�����?=            @U@������������������������       �h{�'@'             N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     Pr@     ��@      8@     �N@     `}@     �V@     Ќ@     `n@     p�@     `u@      @@      @      S@     `e@      @      "@     �X@      ,@     �y@     �H@     �q@     @Q@      @      @      M@      U@               @     �Q@       @     �a@      D@     `a@      G@      @             �G@      R@              @      N@      @     �a@     �@@     �_@      <@      @              D@      J@              @     �D@      @     �]@      6@      X@      4@                      @      4@              �?      3@      �?      5@      &@      >@       @      @      @      &@      (@               @      $@      �?      @      @      *@      2@      �?      @       @      $@               @       @      �?       @       @      $@      2@                      @       @                       @              �?      @      @              �?              2@     �U@      @      �?      =@      @     �p@      "@      b@      7@                      (@     �G@              �?      0@              g@      @     �T@      $@                      @      2@              �?      *@             �\@              J@       @                      @      =@                      @             �Q@      @      ?@       @                      @      D@      @              *@      @     �T@      @      O@      *@                      @     �C@      @              (@      @      I@      @     �G@      *@                       @      �?                      �?             �@@              .@                      6@      k@     �z@      5@      J@     0w@     @S@     �@     @h@     ��@     q@      ;@      $@     �c@     �s@      ,@      @@      o@      N@     `x@      b@     �x@      f@      0@             �M@     �a@      @      @     �U@      "@     �l@     �L@     @i@      P@       @               @     �B@                      3@             �W@      "@      R@      ,@                     �I@      Z@      @      @      Q@      "@     �`@      H@     @`@      I@       @      $@     @X@     `e@      &@      <@     @d@     �I@     @d@      V@     `h@      \@      ,@      @      O@     �Y@      @      0@     �V@      <@     �\@      ?@      ^@      B@      @      @     �A@      Q@      @      (@     �Q@      7@      H@     �L@     �R@      S@       @      (@     �N@     @\@      @      4@     �^@      1@     @^@     �H@     �`@     @X@      &@      (@      M@     �X@      @      2@      [@      0@     �S@      H@      T@     �T@      $@      @      C@     @S@      @      &@     @W@       @     �P@      =@     �P@     �E@      @      @      4@      6@       @      @      .@       @      (@      3@      *@      D@      @              @      ,@               @      ,@      �?      E@      �?     �J@      ,@      �?               @      @                      "@      �?      @@              A@      �?      �?              �?      "@               @      @              $@      �?      3@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJt�%=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @M�� d@�	           ��@       	                    �?����@�           l�@                           �?�1y�	V	@           ��@                           �?�ЄGF@�            �r@������������������������       ��Ih!?@7            @T@������������������������       ���+� @�             k@                            �?Ma��a�	@F           @�@������������������������       �|�=���@�            q@������������������������       �6�t�+�	@�            �n@
                          �5@a�;w~�@|           �@                           �?'���W@�           ��@������������������������       �}����@|            @h@������������������������       �7 $}@6           �~@                            �?/��	@�           ��@������������������������       ��=�Gi�	@�            �w@������������������������       �\�5}�@�            �u@                          �4@�.-��@9           L�@                           @߳���@;           ��@                           @G[2ٙ�?           �z@������������������������       ����G���?�            t@������������������������       �^� @K            �[@                           @�I��@            |@������������������������       ��];��@�            pu@������������������������       �t���@D            �Z@                           @������@�           �@                           �?e��M9@�           `�@������������������������       ��s��@�             y@������������������������       ���q���@�            �w@������������������������       ��#�Z�n@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     �s@      �@      C@     �F@      |@     �S@     ��@      n@     P�@     Pv@      ?@      .@     @n@     �t@      ?@      @@     �r@      M@     `v@      i@     �w@     �n@      >@      @      T@     �^@      5@      (@     �\@      <@     �a@      S@      ^@     @U@      ,@              7@      G@       @       @      E@      @     �S@      4@      I@      4@      �?              @      .@                      ,@              8@      �?      3@      @                      3@      ?@       @       @      <@      @      K@      3@      ?@      0@      �?      @     �L@     @S@      3@      @      R@      5@      O@      L@     �Q@     @P@      *@      �?      5@      H@      @      �?     �A@      .@      =@     �G@     �B@      <@       @      @      B@      =@      0@      @     �B@      @     �@@      "@     �@@     �B@      @      &@     @d@     @j@      $@      4@     �g@      >@     @k@     @_@     pp@     �c@      0@       @      K@     �U@      @      @     �W@      "@     �a@      I@     �c@     �S@      @              4@      8@                      .@             �K@      @      M@      3@               @      A@      O@      @      @     �S@      "@     �U@     �G@     �X@     �M@      @      "@      [@      _@      @      .@     �W@      5@      S@     �R@     �Z@     @T@      $@       @      K@     �K@       @      (@      D@      ,@      B@     �C@     @Q@      F@      @      �?      K@     @Q@       @      @     �K@      @      D@      B@     �B@     �B@      @       @     �R@     �j@      @      *@     `b@      4@     ��@      D@     �z@     @\@      �?             �C@     �Z@      @      @      L@       @     �x@      &@     �k@     �B@                      3@      @@              @      7@             �l@      @      Z@      .@                      3@      2@              @      0@             �f@      �?     �R@      @                              ,@              �?      @              H@      @      =@       @                      4@     �R@      @      �?     �@@       @     �d@      @     �]@      6@                      $@     �J@      �?              5@       @     �a@      @     @W@      .@                      $@      5@      @      �?      (@              7@       @      :@      @               @     �A@     @[@      �?       @     �V@      2@     �l@      =@     �i@      S@      �?       @      @@     @[@               @      U@      .@      l@      9@     `i@      S@      �?       @      7@     @Q@              @      E@      @     @_@       @     �W@      9@                      "@      D@               @      E@       @      Y@      1@      [@     �I@      �?              @              �?              @      @      @      @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJbhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@r�M�aE@�	           ��@       	                    �?��_��i@d           ��@                           @}��I@t           ��@                           �?�r~@           �{@������������������������       �C]�2�@p            �f@������������������������       ��;�I�c@�            pp@                           �?2T�E�@V            ``@������������������������       �`�>�n@              K@������������������������       ���\D6�@6            @S@
                           �?y����@�           ��@                           �?�>}�2 @           @z@������������������������       ����� @�            �l@������������������������       ����S��?t            �g@                          �1@$#+H�=@�           ��@������������������������       �#ZC?�� @�            �o@������������������������       �d�We@E           �@                           @����J@6           Ҡ@                          �<@�^�O��@�           $�@                            @��g��@�           ��@������������������������       �	� k�n@�           �@������������������������       ��dM���@%           �}@                           �?��C�P@�            Pr@������������������������       ���57@G            @]@������������������������       ��,T�@v             f@                            �?�\�P�	@�             l@                          �6@��Ҫ,	@R            �_@������������������������       ��f/��d@             >@������������������������       �s�Fe�@=             X@                           �?Ҭf*P�@;            �X@������������������������       ���<7�F@            �A@������������������������       ���T`P	@#            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     ��@      ;@     �N@     �{@      T@     �@     �h@     ��@     @w@     �B@      @      V@     �l@       @      9@      d@      .@     Ȃ@     �S@     px@     �b@      (@      @      F@     @S@      @      "@     �S@      @     �Y@     �F@      [@      U@      (@       @      ?@      L@       @       @     �J@      @      X@      ?@     �V@      P@      @      �?      @      ;@                      (@      �?      D@      *@      L@      7@              �?      8@      =@       @       @     �D@      @      L@      2@     �A@     �D@      @       @      *@      5@       @      �?      :@       @      @      ,@      1@      4@      @      �?      "@      "@                      "@               @      @       @      *@       @      �?      @      (@       @      �?      1@       @      @      @      .@      @      @              F@     �b@      @      0@     �T@      "@     0@      A@     �q@      P@                      ,@      D@              @      *@              l@      @     @X@      2@                      $@      3@              @      $@             �_@      @     �E@      "@                      @      5@                      @             @X@       @      K@      "@                      >@     �[@      @      "@     @Q@      "@     0q@      ;@     @g@      G@                      @     �B@              �?      &@             �[@      &@     �Q@       @                      ;@     �R@      @       @      M@      "@     �d@      0@     �\@      C@              $@      j@     �u@      3@      B@     �q@     @P@     �x@     �]@     �z@      l@      9@      @     `f@     �s@      1@     �A@      o@      J@     �v@     �U@     @y@      j@      .@      @     �b@     �p@      0@      ;@     @j@      E@      u@      P@      v@      c@      (@      @      X@     @h@      @      7@     �a@      C@      n@      @@     �p@     �Z@       @             �K@     �Q@      "@      @     �Q@      @     �W@      @@     @V@      G@      @              <@      H@      �?       @     �C@      $@      ;@      7@      I@      L@      @              @      >@              @      "@       @      (@      @      4@      5@                      7@      2@      �?      @      >@       @      .@      0@      >@     �A@      @      @      >@      A@       @      �?     �@@      *@      >@      ?@      5@      0@      $@      �?      5@      .@       @      �?      $@      &@      .@      :@      ,@      @      @              @      @      �?      �?      @      @      @      �?              @              �?      0@      "@      �?              @      @      &@      9@      ,@      @      @       @      "@      3@                      7@       @      .@      @      @      "@      @       @      �?      @                      @       @      @       @      �?      "@      �?               @      .@                      0@              "@      @      @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��J`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?&��/@�	           ��@       	                    �?LW�  @&           �@                           �?Ś8&�t@�           0�@                          �;@�A��,�@�             k@������������������������       �q.aG�@x             g@������������������������       ��8�Rj@             @@                            �?
}P�@'           �|@������������������������       ��ѕ�>5�?H            �\@������������������������       ��[IW�@�            �u@
                           �?��>&�@r           ؂@                          �<@Dv-4"�@�            p@������������������������       �5����\@�            �l@������������������������       �ts �� @             ;@                           @���}�i@�            �u@������������������������       ���h@>             Z@������������������������       �c���K@�            @n@                            @�m�L)@�           ��@                           @O��n��@�           ��@                           @@���a!	@;           (�@������������������������       �X@����@&            �@������������������������       ��-ZmZ@            �@@                          �6@C����7@]           Ѝ@������������������������       �i���2@�           ��@������������������������       ����#:@�            �r@                           �?s�	 	@�           H�@                           @#i��	@?           �@������������������������       �f�W�T	@�             u@������������������������       �#�x	@h            �e@                           �?M��#W@�            �p@������������������������       ��%�K�@H            �Y@������������������������       �\�md@�@o            `d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@      s@     Ё@      @@     �K@      |@      N@     0�@     @j@     ��@     �v@     �C@             �S@      g@      �?      @     @]@      "@     �}@      E@     �q@     �S@      @              C@      W@      �?      @      M@      @     �q@      7@     ``@      C@      �?              5@      @@      �?      @      =@      �?     �K@      .@      B@      6@      �?              5@      ;@      �?       @      7@              K@      $@      ?@      ,@      �?                      @              �?      @      �?      �?      @      @       @                      1@      N@              @      =@       @      m@       @     �W@      0@                              $@              �?      "@      �?     @P@              9@      @                      1@      I@               @      4@      �?     �d@       @     �Q@      (@                      D@     @W@              �?     �M@      @     `g@      3@     @c@      D@      @              9@     �H@              �?     �D@              F@      &@     �M@      9@       @              7@     �F@              �?     �B@             �E@      $@      M@      &@       @               @      @                      @              �?      �?      �?      ,@                      .@      F@                      2@      @     �a@       @     �W@      .@       @              @      @                      @      @      B@      �?     �E@      @                       @     �C@                      ,@       @     �Z@      @      J@      &@       @      $@     @l@     x@      ?@      H@     �t@     �I@     ��@      e@     `@     �q@      A@       @     �a@     p@      3@      B@      l@     �@@      {@     �]@      w@     �i@      .@      �?     �U@     �`@      *@      ;@     �^@      7@     �a@      W@      `@     �^@      *@              T@     @`@      *@      ;@     @]@      6@     �a@      V@     �^@      ^@       @      �?      @       @                      @      �?              @      @       @      @      �?      L@     @_@      @      "@     �Y@      $@     `r@      ;@     �m@     �T@       @              :@     �U@      @       @      Q@      @      n@       @     �b@      L@       @      �?      >@     �C@       @      �?      A@      @      K@      3@      V@      ;@               @      U@      `@      (@      (@     �Z@      2@      `@     �H@     �`@     �S@      3@       @     @Q@     �R@       @      @     �S@      .@     @P@     �D@     @S@     �I@      3@       @     �G@     �I@       @      �?     �L@       @     �E@      9@     �I@      >@      "@              6@      7@              @      5@      @      6@      0@      :@      5@      $@              .@      K@      @      @      <@      @     �O@       @     �L@      <@                       @      2@      @      �?      $@      @      6@      @      =@      (@                      *@      B@      �?      @      2@             �D@      @      <@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�NOhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@��@�	           ��@       	                    �?�Kԇ"J@}           ��@                           @,oC��i@�           �@                          �1@���G@�            �r@������������������������       �3:� @8             X@������������������������       ��i�9@�             i@                          �0@��=�q< @�            �w@������������������������       �\Q��T�?"            �I@������������������������       �4��3� @�            �t@
                           @%��0/�@�           ��@                          �2@B*\�*@�           8�@������������������������       ��ZK'[]@e           0�@������������������������       ��`���}@(           �|@                           @�p6M۵@J            @\@������������������������       �7g�B�	@+             O@������������������������       ��<ު��@            �I@                           �?�D�]u�@?           N�@                          �<@?̥a�r@f           X�@                           @w�;��@-           �}@������������������������       ��#/�p�@�             r@������������������������       ���Uxj�@q            �f@                            �?�*�_a�@9            �T@������������������������       �m�*���@             6@������������������������       ��Sv3J�@-            �N@                          �:@�|���;	@�           �@                          �5@Ǟ�� �@�           ܐ@������������������������       �0��]��@�            �k@������������������������       ��C���@(           Ȋ@                           @�J�*=	@           P|@������������������������       ���HRE	@�            ps@������������������������       ���5䵳@V            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     ؀@      5@     �P@      |@     @W@     H�@     �k@     @�@     �w@      =@      @     @X@     `m@      @      5@     `f@      1@     ��@     @U@     �y@     �`@      $@              B@     �R@               @      L@      �?     `r@      4@     `c@     �B@                      2@      C@                     �A@      �?     �V@      .@     @S@      5@                      �?      &@                      ,@              D@      @      :@      �?                      1@      ;@                      5@      �?     �I@      (@     �I@      4@                      2@      B@               @      5@             `i@      @     �S@      0@                              (@                      @              <@               @      @                      2@      8@               @      .@             �e@      @      S@      *@              @     �N@      d@      @      3@     �^@      0@     �t@     @P@      p@      X@      $@      @      L@     �b@      @      0@     @[@      *@     0s@     �J@     `n@      S@      @      �?      =@     @Y@      @      �?     @P@      �?     �g@      ;@     ``@     �@@              @      ;@     �H@       @      .@      F@      (@     @]@      :@      \@     �E@      @      �?      @      &@              @      ,@      @      9@      (@      *@      4@      @      �?      @      @              @      (@      @      @      $@      "@      @      @               @      @                       @              6@       @      @      *@              ,@      k@      s@      0@      G@     �p@      S@     pu@     @a@     �x@     �n@      3@             �G@     @V@       @      @      F@      "@     `a@      :@      `@      N@      @             �D@      T@       @      @      ?@      "@     @`@      4@      \@     �D@      @              B@      E@       @      @      :@       @     �P@      ,@     @P@      ?@      @              @      C@                      @      @      P@      @     �G@      $@                      @      "@              @      *@              "@      @      1@      3@      �?              @      @                      @                       @      @      �?      �?               @      @              @      @              "@      @      *@      2@              ,@     @e@     �j@      ,@      D@     `l@     �P@     �i@      \@     �p@     @g@      .@      @     �[@     �e@      $@      ;@      e@     �H@     �d@      S@     �g@     @W@      *@       @      @     �E@      �?      @      E@      *@      6@      *@     �J@      0@      @      �?      Z@     ``@      "@      4@     �_@      B@     �a@     �O@      a@     @S@      $@      &@     �M@     �D@      @      *@      M@      2@      D@      B@     �S@     @W@       @      &@      B@      ?@      @      "@      ;@      2@      3@      A@      F@     @S@       @              7@      $@      �?      @      ?@              5@       @      A@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�PlEhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @E�l��'@�	           ��@       	                   �<@< ��@�           6�@                           �?d���Q@�           ��@                           �?���@�           �@������������������������       ����l}�@            {@������������������������       ���doT	@v           ��@                           �?1ۜ&�6@[           �@������������������������       �!n���@�             l@������������������������       ��B�@�            �s@
                           �?/QF	@�            `o@                           �?����@:            @T@������������������������       ���LЬ1@
             .@������������������������       ��lҔ��@0            �P@                          �@@s�b�ct	@f            @e@������������������������       �w�n��@[             c@������������������������       ��F:�@             2@                          �1@qJ�q�@2           ��@                           @j�Q�B�?�            �t@                            �?�!����?�            �o@������������������������       �I�w�"�?\            �a@������������������������       ��SjI�?L             \@                           @~g<�=�@2            @S@������������������������       �a��@(             O@������������������������       �E��I�d�?
             .@                           @3��V�@X           ��@                          �:@���.��@D           x�@������������������������       �����D�@            �@������������������������       �7P�4�3@?            �Z@                           �?�+��6:@           @{@������������������������       �Ӫ5@Vl@a             c@������������������������       �8r2ph@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     @q@     (�@     �@@     �J@      ~@     @R@     X�@     �j@     P�@     �v@      <@      1@     �h@     �t@      5@      B@     �t@     �L@     Px@      g@     v@     0p@      9@      *@     �e@     �r@      1@      <@     �r@      D@     `w@     �b@     �t@     �h@      7@      *@     �`@     @l@      1@      6@     �l@      ;@     @l@     �\@     �k@     �c@      7@      �?      C@     �Q@      @      @      O@       @     �Y@      5@      V@      A@      @      (@     @X@     `c@      ,@      2@      e@      9@     �^@     @W@     �`@     �^@      2@              C@     @S@              @      Q@      *@     �b@      B@     @\@      E@                      @      ?@               @      A@      "@     @P@      ,@      E@      4@                      ?@      G@              @      A@      @     �T@      6@     �Q@      6@              @      9@      @@      @       @      ?@      1@      .@      A@      3@      N@       @      �?      "@      (@              @      &@               @      (@      @      7@      �?              @      @                       @                              �?      @              �?      @      "@              @      "@               @      (@      @      3@      �?      @      0@      4@      @       @      4@      1@      *@      6@      .@     �B@      �?              ,@      3@      @       @      1@      ,@      (@      6@      .@     �@@      �?      @       @      �?      �?              @      @      �?                      @                     �S@     �j@      (@      1@     �b@      0@     ��@      ?@     �z@     �Z@      @               @     �D@              @      "@             �g@             �R@      *@                       @      <@                      @              d@              J@      @                      �?      &@                       @             @X@              8@      @                      �?      1@                      @             �O@              <@                                      *@              @      @              <@              6@      @                              *@               @      @              7@              ,@      @                                               @                      @               @                              S@     �e@      (@      *@     �a@      0@     P}@      ?@     �u@     @W@      @              I@     �\@      @      @     �W@      "@     `u@      .@     �n@      O@       @              F@     �X@      @      @     �Q@      "@      t@      .@     �j@     �J@       @              @      0@                      8@              4@              @@      "@                      :@     �M@       @      "@      H@      @     �_@      0@      Z@      ?@      �?               @      6@       @      �?       @      @     �P@      @      @@      @                      2@     �B@      @       @      D@      @     �N@      &@      R@      9@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�+q<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��s�Vo@�	           ��@       	                    �?uī�@�           ,�@                           �?�
s�@'           �~@                            �?0BQȍw@            `k@������������������������       �!?��j�@?            @]@������������������������       �p,��N~@@            �Y@                           �?{-D��@�            q@������������������������       ����4�@E             ]@������������������������       �s�O���@c            �c@
                            �?��%	0@�           ��@                           @$���S@r            `h@������������������������       �ۿI2yf@(            @P@������������������������       �X�0#>@ @J            @`@                            @u�L���@V           ��@������������������������       ��+/+�@           �y@������������������������       ��r��K* @T             `@                           @;x���S@�           ��@                           �?��)@�           p�@                           @>Ɂ{�	@p            �f@������������������������       �u+��@L             `@������������������������       �{�4K��@$             J@                           �?�+ l�@           �@������������������������       �X�{�]�	@�           ��@������������������������       ��X;U@u           ��@                          �5@���4H@2            �Q@                            �?�Y�Sv@             =@������������������������       �|R��>@             0@������������������������       ����aM@             *@                           �?��Ef�@            �D@������������������������       �����Z@             "@������������������������       �͠&Ί@             @@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     Pu@     P�@      A@     �O@      |@     @R@     ��@      k@     ��@     `w@      >@             @Y@     @d@      @      @     �X@      (@     P{@     �F@      q@      U@      @              N@     �R@      @      @      L@      �?     @[@      A@      X@      J@      @              3@      ;@      @      @      <@      �?     �G@      4@      F@      9@      �?              ,@      0@       @       @      $@              9@      $@      3@      2@      �?              @      &@       @      �?      2@      �?      6@      $@      9@      @                     �D@     �G@                      <@              O@      ,@      J@      ;@       @              .@      3@                       @              :@      @     �@@      "@       @              :@      <@                      4@              B@      $@      3@      2@                     �D@      V@              �?      E@      &@     �t@      &@     @f@      @@      @              @      1@              �?      *@      "@      W@      @     �F@      "@       @              @      @              �?      @      @      3@              9@       @       @                      &@                      $@      @     @R@      @      4@      @                      C@     �Q@                      =@       @     �m@      @     �`@      7@      �?              ?@     �O@                      4@       @     �e@      @     �X@      1@      �?              @       @                      "@             �O@      �?     �A@      @              0@      n@     �x@      >@     �M@     �u@     �N@     ��@     `e@     �}@      r@      8@      *@     �l@     @x@      =@     �M@     u@      L@     ��@     �c@     p}@     �q@      5@              >@      2@              "@      ;@      "@      2@      7@      9@      4@       @              ;@      (@              "@      8@       @      @      .@      $@      1@       @              @      @                      @      �?      *@       @      .@      @              *@     �h@      w@      =@      I@     `s@     �G@     `�@     �`@     �{@     `p@      3@      *@     �\@      e@      5@     �@@     �d@     �B@     �_@     �U@      `@     �b@      .@              U@     @i@       @      1@      b@      $@     �z@     �G@     �s@     �\@      @      @      &@      @      �?              *@      @              ,@       @       @      @       @       @      �?                      @      @                      @      @       @      �?       @                                       @                      @      @      �?      �?              �?                      @       @                              @      �?      �?      "@      @      �?               @      �?              ,@       @      �?      �?      �?                                      @                       @      �?      �?      �?              "@      @      �?              @      �?              (@      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��MVhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�a���@�	           ��@       	                    �?d���&�@u           ��@                          �<@��.�z@�           �@                           �?![<��@e           (�@������������������������       ��XUh�?@�            pq@������������������������       �%�h�2�@�            �r@                           �?�̇�'9@*             N@������������������������       ��"-��@             <@������������������������       �t(#�]�@             @@
                          �3@��+Q	@�           <�@                            �?L�0���@0           p~@������������������������       �5�5�fd@\            `b@������������������������       ���hj�@�            @u@                           �?m���t�	@�           ��@������������������������       ����:�	@           (�@������������������������       ���-���@�            0r@                           �?�	�%�@1           �@                            @���9@c           ��@                          �5@:a�A�@            {@������������������������       �sfX�X @�            �r@������������������������       ���{���@P            @`@                          �2@F�w�K�?D             [@������������������������       �u�C�$ �?              J@������������������������       ��'U��� @$             L@                           �?�-�w��@�           t�@                           @Dep��;@P           �@������������������������       ������E@�            `w@������������������������       ����*Y�@Z            �a@                          �7@^���@~           ؂@������������������������       �VQs�fh@           `{@������������������������       �a�).��@l            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     X�@     �@@     �J@     �|@     �T@     @�@     @m@     ��@     0x@      A@      ,@     �j@     Pv@      5@     �E@     Pt@     @P@     �v@     �g@     0x@     �o@      <@      �?     @P@      W@      @      @      Q@      @     �c@      B@      c@      J@      @      �?      N@     �T@      @      @     �M@      @     �c@      :@     `b@     �A@       @      �?      >@     �A@      @      @      @@      @     @R@      4@      M@      0@       @              >@      H@                      ;@             �T@      @     @V@      3@                      @      "@              @      "@              �?      $@      @      1@      �?              �?      @              �?       @                      @       @      *@                      @      @               @      @              �?      @      @      @      �?      *@     �b@     �p@      2@     �B@     p@     �M@     `i@      c@     `m@      i@      9@       @      B@      S@      �?      �?     �N@      "@      W@      H@     @S@     �R@      "@              ,@      5@                      7@      �?      =@      1@      8@      (@      @       @      6@     �K@      �?      �?      C@       @     �O@      ?@     �J@     �O@      @      &@     @\@     �g@      1@      B@     �h@      I@     �[@     @Z@     �c@     �_@      0@      &@     �T@      a@      .@      =@     �a@     �C@     @Q@     �V@     �[@      Y@      .@              >@     �J@       @      @      L@      &@      E@      .@      H@      :@      �?             @V@     �l@      (@      $@     �`@      2@      �@     �F@      y@     �`@      @              7@     �S@               @      8@      @     �o@       @     �_@      6@                      2@      S@              �?      4@      @      h@      @      X@      3@                      (@      H@              �?      .@       @      d@      @      J@      @                      @      <@                      @      �?     �@@      �?      F@      (@                      @      @              �?      @             �M@       @      ?@      @                       @      �?                                      B@              &@       @                      @       @              �?      @              7@       @      4@      �?                     �P@     �b@      (@       @     �[@      .@     @t@     �B@     0q@      \@      @              E@      P@      @      @     �O@      @     �_@      .@     @`@      K@      @              =@     �G@              �?      G@      �?     �[@      (@     �U@     �B@      @              *@      1@      @      @      1@       @      1@      @      F@      1@                      8@     �U@      @      @      H@      (@     �h@      6@      b@      M@      �?              2@      S@      @      �?      5@      @      e@      @     �Y@      @@      �?              @      &@       @       @      ;@      @      <@      .@     �E@      :@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���LhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��A��U@�	           ��@       	                    �?,� #	@�           ��@                          �<@nT ǋ�@-           �~@                           �?ϼ�<�@           �{@������������������������       �h/�h�@h            �d@������������������������       �5s֊�<@�            pq@                          �>@[���U@"             H@������������������������       �h}�X��?             6@������������������������       �}�6@             :@
                           �?�s.ñ	@�           �@                            �?�D�c��@           0{@������������������������       �\@'	�E@W             `@������������������������       ���lV��@�             s@                            �?.��"�Q
@�           8�@������������������������       �1_�Y
@�             v@������������������������       ������	@�            pv@                           �?�Vp�>@�           ȡ@                          �7@S�Z�@�           p�@                          �4@p�"�@z           ��@������������������������       �I#�I���?            |@������������������������       �$����@\            �b@                           @@�1��W�@_             c@������������������������       �T+�n@X            `a@������������������������       �rD��*@             ,@                          �4@�7�7Gs@�           ؗ@                            �?�H݇�@�           �@������������������������       �ro�*�@	           @z@������������������������       ��>
���@�            �s@                           @:�W*�@�           ��@������������������������       �����i@�           ��@������������������������       �9//"�@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     @q@     X�@      @@     �O@     �{@     �T@      �@     �k@     (�@     0x@      ;@      2@     `b@     �o@      7@      B@     `l@     �E@     0p@     �`@     �o@     �k@      3@             �H@     @R@      @      @     �N@      @     �^@      6@     @X@     �I@      @              G@      Q@      @       @      K@      @     �]@      1@     �W@      ?@      @              "@      7@                      9@              K@      @      E@       @                     �B@     �F@      @       @      =@      @     @P@      ,@     �J@      7@      @              @      @               @      @              @      @       @      4@                      �?      @                                      �?      �?              .@                       @      �?               @      @              @      @       @      @              2@     �X@     �f@      2@      @@     �d@      D@      a@     @\@     �c@     �e@      0@       @      5@     �S@      @       @      N@       @     �S@     �C@      M@      S@       @              @      *@              @      5@      @      =@      *@      7@      2@      �?       @      1@     �P@      @      @     �C@      @     �H@      :@     �A@      M@      �?      0@     @S@     �Y@      ,@      8@     �Z@      @@      M@     �R@     �X@      X@      ,@      @      G@     �H@      @      .@      C@      .@      9@     �G@      D@     �K@      $@      "@      ?@     �J@      "@      "@      Q@      1@     �@@      ;@      M@     �D@      @      �?      `@     �r@      "@      ;@     @k@     �C@     (�@     �U@     @�@     �d@       @             �@@     �T@       @       @      E@       @     �u@      *@     `g@     �@@       @              >@     �Q@       @       @     �B@      @     pr@      @     �`@      1@       @              5@      D@               @      6@             `m@      @     �[@      (@       @              "@      ?@       @              .@      @      N@              8@      @                      @      (@                      @      @      I@      "@     �J@      0@                      �?      (@                      @       @      I@      @     �I@      (@                       @                                      @              @       @      @              �?      X@     @k@      @      9@      f@      ?@     �z@     �R@     �t@     ``@      @             �B@      Z@      @       @     �L@      @     `p@      ?@     �d@      O@                      2@     �H@       @      @      A@      �?     @b@       @     �[@     �F@                      3@     �K@       @       @      7@      @      ]@      7@      L@      1@              �?     �M@     �\@      @      1@     �]@      8@     �d@     �E@     �d@     @Q@      @      �?      L@     @\@       @      1@      [@      6@     �d@      B@     `d@      Q@      @              @      �?      �?              &@       @              @      @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�L0;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�u�p4b@~	           ��@       	                     @&B��@�           ��@                           @y$\�@)           Ћ@                           �?�vJ��@	            {@������������������������       ���5�s�@~            �i@������������������������       ���E*C,@�            �l@                           @f�z�o@            �|@������������������������       ��$hW^�?�            �s@������������������������       ����'@_            �a@
                           �?��⻽�@�            Pt@                          �8@�cd��@m            @g@������������������������       ��E���@P             `@������������������������       �8a�Sm�@             M@                           �?2]�T8^@W            `a@������������������������       �/K��@8             V@������������������������       ��H��?            �I@                          �7@���0e&@�           �@                           @aI�|�I@x           p�@                          �1@�4E��6@�           @�@������������������������       �ٽ��F@�            @k@������������������������       ���$`��@U           ��@                          �3@���@�           `�@������������������������       ����d��@�            s@������������������������       �8r~�@�            �u@                          �:@�z��
	@           p�@                           �?Z	Gh�@           pz@������������������������       �Ulѣ@            �@@������������������������       ���A��@�            `x@                           @"�QIb�@           p|@������������������������       �e
��f@{            @k@������������������������       ��d�g@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     0�@      >@     �I@     @}@     �T@     `�@      n@      �@     pw@      ?@      �?     @S@     @e@      @      &@     `a@      (@     p{@      K@     �l@     �R@      @      �?      F@      b@      @      @     @W@      (@      t@      ?@      f@      K@      @      �?     �@@     �L@       @      @     �P@      @     �Z@      9@     �V@     �B@      @      �?      @      :@       @      @     �A@      @      G@      .@      C@      8@      @              :@      ?@              �?      @@      �?     �N@      $@     �J@      *@                      &@     �U@       @      �?      :@      @     �j@      @     @U@      1@                      @      M@                      3@      @     �d@       @     �I@      @                      @      =@       @      �?      @      @      H@      @      A@      $@                     �@@      :@      �?      @      G@             @]@      7@      K@      4@                      6@       @      �?      @      9@              Q@      ,@      @@      &@                      &@      @      �?              (@              L@      @      9@      "@                      &@      �?              @      *@              (@      @      @       @                      &@      2@                      5@             �H@      "@      6@      "@                      &@      0@                      2@              7@      @      @      "@                               @                      @              :@      @      1@                      *@     `k@     �y@      9@      D@     �t@     �Q@     ��@     @g@     �@     �r@      <@      @      `@     �r@      .@      ?@     �j@      D@     �|@     �U@     v@      e@      *@      @     �Q@      g@      ,@      0@      b@      ?@     �q@      L@     �o@     �[@      @               @      <@                      ,@             @Q@      ,@     �P@      2@              @      O@     �c@      ,@      0@     @`@      ?@     �j@      E@      g@      W@      @       @      M@     �]@      �?      .@     @Q@      "@     �f@      ?@     @Y@     �M@      "@              6@     �D@              @      5@      @      [@      .@      H@     �B@      @       @      B@     @S@      �?      &@      H@      @      R@      0@     �J@      6@      @      @     �V@     @[@      $@      "@      ]@      >@      Z@     �X@     �c@     �`@      .@             �C@     �K@      @      @      M@      1@      J@      H@     @V@      G@      $@              @      @               @      "@              �?      @      @       @                      @@      J@      @      @     �H@      1@     �I@      E@     �U@      F@      $@      @      J@      K@      @      @      M@      *@      J@     �I@      Q@     �U@      @      @      0@      B@      �?      @      >@      @      4@      <@      1@     �J@      @       @      B@      2@      @      �?      <@      @      @@      7@     �I@     �@@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJr4�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @x�.3�?@�	           ��@       	                    �?���)�@j           F�@                           �?���"o>	@�           H�@                          �<@�;��Z@#           �|@������������������������       �/d.nէ@            0y@������������������������       �N-�W�@#            �L@                          �4@8~���	@�           �@������������������������       �w�φd@�             z@������������������������       ������	@�           0�@
                            �?�QΥ�@�           ��@                           �?"Ն��@�             u@������������������������       �L*��o@Z             a@������������������������       �'z���@~            @i@                          �4@���E7@�            �o@������������������������       �+��k�J@M             ^@������������������������       �Id�U@[            �`@                           �?ױ�I��@3           ��@                           @�oE�/@v           ��@                          �2@g5�N:��?�            Px@������������������������       ����<D�?r            `f@������������������������       �/�w@�            @j@                          �5@8$Qf��@�             j@������������������������       ����^<@Z            �a@������������������������       �c6K��@*            @Q@                          �<@"�`;��@�           @�@                           @Ðp��@�           H�@������������������������       �~��x.@�           ȏ@������������������������       ��E��@             9@                           @�>�(�$@(             O@������������������������       �9�)��r@             A@������������������������       �ɖnL(��?             <@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     0r@     ��@      ?@      G@      }@     �T@     �@     �k@     ��@     0x@      :@      1@      j@     Pt@      7@      C@     0u@     �N@      w@      f@     Pw@     p@      9@      1@     �b@     �l@      5@     �@@     @p@      J@      n@      a@      o@     �i@      6@              >@     �Q@      �?      "@     �N@             �\@      <@     �W@     �H@      @              ;@      Q@      �?      @      K@             �[@      5@     �U@      ;@      @              @      @              @      @              @      @       @      6@              1@     @^@      d@      4@      8@     �h@      J@     �_@      [@     `c@     �c@      3@       @     �B@      E@      $@      @     �Q@      "@      S@      >@     @S@      K@      @      .@      U@     �]@      $@      4@      `@     �E@      I@     �S@     �S@     �Y@      .@             �L@     �W@       @      @     �S@      "@      `@     �D@      _@     �I@      @             �A@     �D@       @      @      C@      @     �P@      3@      W@     �@@      @              .@      5@               @      3@      @      =@      $@      8@      (@      �?              4@      4@       @      �?      3@      @     �B@      "@      Q@      5@       @              6@     �J@               @     �D@      @      O@      6@      @@      2@                              :@               @      4@      �?     �B@      *@      ,@      @                      6@      ;@                      5@       @      9@      "@      2@      &@                     �T@     @j@       @       @     �_@      6@     h�@      F@      |@     @`@      �?              4@     �S@      @              2@      @     0r@      *@      a@      ?@                      .@      H@                       @      @     �i@      @     �U@      0@                      @      1@                      �?             �]@              A@      @                      $@      ?@                      @      @     �U@      @     �J@      *@                      @      ?@      @              $@             �U@      $@     �H@      .@                      @      7@                      @             �P@      @      <@      @                               @      @              @              4@      @      5@       @                     �O@     ``@      @       @     @[@      .@     �t@      ?@     �s@     �X@      �?              L@     @_@      @      @     @V@      .@      t@      ?@     �r@      W@      �?              K@     @_@      @      @     @U@       @     t@      >@     �r@      V@      �?               @                       @      @      @      �?      �?      @      @                      @      @      �?       @      4@               @              &@      @                      @      @      �?       @      @              @              @      @                      @                              *@              �?              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��j{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�Mn��1@�	           ��@       	                    �?��5s�@�           p�@                           �?�ꢊ�"@&           �}@                           �?�(s4�<@n            �e@������������������������       ���PS�@6            @S@������������������������       ��im�o	@8            �W@                           �?�@X�j@�            �r@������������������������       ��$��*1@W            �a@������������������������       ��	Ʃ�@a            �c@
                            @���6�@�            �@                          �=@�ia3.@s           (�@������������������������       ��T�I<�@g           ��@������������������������       ��(;��e@             3@                           7@6Hs�?Y            �c@������������������������       ��e�i� �?F            @`@������������������������       ������,�?             =@                           @�>�@�           ڤ@                          �5@��A��n	@�           ��@                           �?�|���@�           0�@������������������������       ���K�}@�             n@������������������������       �<�wB@.           `}@                          �6@�n6�
@           ȉ@������������������������       �\�w�V@Z             b@������������������������       �>U#
@�           @�@                           �?J�~Q��@�           ��@                           @�7�V@b           ��@������������������������       ��֕�@@           �~@������������������������       ����jeK@"            @P@                           @9��{�3@e           ��@������������������������       ��H�#S@�            py@������������������������       ����Ks$@k            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     0s@     ��@      @@     �J@      {@     �R@     T�@     �j@     Ј@     �u@      @@       @     �V@      f@      @      "@     �Z@      "@     �{@      A@     `q@     �U@      @       @      L@     �S@      �?      @     �N@      @     �V@      2@     �W@     �L@      @       @      5@      1@                      0@              I@      @     �B@      8@      �?       @      "@      @                       @              7@       @      2@      &@                      (@      *@                       @              ;@       @      3@      *@      �?             �A@     �N@      �?      @     �F@      @      D@      ,@      M@     �@@       @              &@      5@      �?      @      8@      @      7@      $@      7@      3@                      8@      D@              �?      5@              1@      @     �A@      ,@       @              A@     �X@       @       @     �F@      @     0v@      0@     �f@      >@       @             �@@      V@       @              A@      @     �p@      ,@     �a@      5@       @              @@      V@       @              @@      @     �p@      $@     �a@      .@                      �?                               @              �?      @      @      @       @              �?      $@               @      &@              U@       @      D@      "@                              "@               @      &@             �P@              B@      @                      �?      �?                                      2@       @      @      @              0@      k@     x@      =@      F@     �t@     �P@     ��@     @f@      �@     pp@      ;@      ,@      c@     `m@      7@      A@     �m@      J@     @k@     �b@     `l@     `e@      7@      @      H@     �Y@      @      *@     �^@      (@     �b@      L@     �^@     �P@      @       @      2@     �D@      @      @     �G@      @      D@      6@      ;@      <@       @       @      >@      O@       @      $@      S@      @     �[@      A@     �W@     �C@      @      $@     @Z@     �`@      2@      5@     @\@      D@     �P@     @W@     @Z@      Z@      1@      �?      :@      5@              @      1@      @      1@      6@      5@      "@              "@     �S@     �[@      2@      ,@      X@      B@      I@     �Q@      U@     �W@      1@       @      P@     �b@      @      $@      W@      ,@     �w@      =@     r@      W@      @       @      C@     �T@      �?      "@     �G@       @     �e@      1@     �b@     �C@      @       @      9@     �R@      �?      @      F@              d@      &@      a@     �A@      �?              *@      @              @      @       @      (@      @      (@      @       @              :@      Q@      @      �?     �F@      (@     @j@      (@     �a@     �J@      �?              $@      J@      �?              ?@      @     �d@       @     �Z@      >@                      0@      0@      @      �?      ,@      "@     �F@      @      A@      7@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ҃�2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?;�Mgd@�	           ��@       	                    �?��ڒ�@           ȓ@                           �?�?��k@9           @                          �8@����'@�            �k@������������������������       ��M�w��@b            �b@������������������������       ���^	@+            �R@                            @Y{�g�@�             q@������������������������       �#܆�|P@p             e@������������������������       ��y���_@<            @Z@
                           @z�Z�	@�           �@                            �?mԆ�[Q@U           P�@������������������������       ����H�?P            @_@������������������������       ��`%�t�@           �z@                          �5@���B\@�            �j@������������������������       ��ֵ~'�@N            �_@������������������������       �ȏ���U@7             V@                           �?�z��:@�           ��@                           �?L�t@a�	@�           0�@                            �?n�&[�@�            �x@������������������������       �/���@L             ^@������������������������       ��N@�d@�            `q@                           �?��n���	@�           ��@������������������������       �+Dw�~	@�            �l@������������������������       �s$���	@(           p}@                           @F�q��V@�           ,�@                            �?7=���@           �{@������������������������       �P^���@V            `a@������������������������       �i�5GdQ@�            �r@                          �5@�,��4�@�           D�@������������������������       �Mb��ב@�           0�@������������������������       �I2	�@           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �u@     X�@      7@      M@     �{@     @T@      �@     `j@     ��@     pu@     �C@              Z@     �d@      @      1@      Y@      &@     p{@     �C@     �r@     �R@      @             �Q@     �Q@      @      (@      H@      @     �X@      <@      [@     �H@      @              <@      4@      @      @      6@      @     �I@      7@     �F@      1@      @              ,@      *@      @       @      ,@      �?      G@      ,@      @@      @      @              ,@      @              @       @       @      @      "@      *@      (@                      E@     �I@              @      :@              H@      @     �O@      @@       @              5@      ?@               @      6@              5@      �?      H@      5@       @              5@      4@              @      @              ;@      @      .@      &@                      A@      X@      �?      @      J@       @     @u@      &@     @h@      :@       @              =@     @Q@              �?      A@      @      p@      "@     �`@      *@                       @      3@              �?      @      �?     @P@              >@      @                      ;@      I@                      >@      @      h@      "@     @Z@      $@                      @      ;@      �?      @      2@       @     �T@       @     �M@      *@       @              @      3@              @      @              L@      �?      ;@      @       @                       @      �?              (@       @      :@      �?      @@      @              0@     �n@     @z@      2@     �D@     �u@     �Q@     h�@     �e@      }@     �p@      @@      0@     @]@     �e@      ,@      7@     �d@      G@     �`@     @[@     �a@     `b@      2@      �?      >@     �P@       @      .@      P@      $@     @P@      >@      M@     �J@      @              (@      *@              @      4@      @      5@      ,@      7@       @              �?      2@     �J@       @      &@      F@      @      F@      0@     �A@     �F@      @      .@     �U@     �Z@      (@       @      Y@      B@     �P@     �S@     �T@     �W@      ,@       @      7@     �G@      "@      @      4@      $@      .@      @@      :@      E@       @      *@      P@      N@      @      @      T@      :@      J@     �G@     �L@      J@      (@              `@     �n@      @      2@     �f@      8@     �z@     �O@     0t@     @^@      ,@             �G@     �Q@      �?      @      M@      (@     @X@      A@     �Q@     �F@      �?              @      9@               @      .@      @      C@      @      3@      5@      �?              E@      G@      �?      @     �E@      @     �M@      <@     �I@      8@                     @T@      f@      @      (@     �^@      (@     �t@      =@     �o@      S@      *@              A@     �]@      �?       @      K@      @      l@      (@      e@      D@      (@             �G@     �L@       @      @      Q@      @      Z@      1@     @U@      B@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO NhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��Q�U�@�	           ��@       	                   �1@c\=B��@j           �@                           �?m�DX�@�           8�@                          �0@�5k�4�@�            r@������������������������       �#��N�@<            �W@������������������������       ��g�y� @�            @h@                           @Xx�*+@�            `t@������������������������       �L�n=$B@g            @d@������������������������       �$���k�?c            �d@
                           �?�&����@�           ��@                           @X�b�a�@2            �@������������������������       ��U����@�            �s@������������������������       ����or�?o            �h@                           @��S*��@�           ��@������������������������       ��4"e^	@t           Ё@������������������������       �W���ǳ@=           �~@                           �??��{��@8           �@                          �>@�D�E@           P{@                            �?��,��@�             x@������������������������       �֑�T'i@F            @\@������������������������       �Po��P@�            q@                          �@@x��=@            �I@������������������������       �l����v@            �@@������������������������       ��xe�_@
             2@                          �?@e��[s	@(           �@                           @6C��:	@�           ��@������������������������       �;�|��	@�           ؇@������������������������       ��!G�|�@           �z@                            �?���0Y�	@:            @W@������������������������       ���s��@             G@������������������������       �[�Ay��@            �G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@      t@     ��@      9@      K@     p{@     �Y@     �@     �j@      �@     �u@     �@@      $@     �^@     pt@       @      7@      j@     �F@     ��@     �U@     @~@     �e@      (@      �?      8@     �W@      �?      �?     �C@       @     �o@      3@     @b@     �A@              �?      "@     �F@      �?              2@       @      `@      "@     �I@      9@                      �?      1@                       @              D@       @      4@      @              �?       @      <@      �?              $@       @      V@      @      ?@      2@                      .@      I@              �?      5@              _@      $@     �W@      $@                      (@      =@              �?      2@              G@      @      E@      @                      @      5@                      @             �S@      @     �J@      @              "@     �X@      m@      @      6@     @e@     �E@     p{@     �P@      u@     `a@      (@              ?@     �S@               @      B@      @     �h@      1@     �\@     �@@                      9@      I@                      <@      @     @W@      1@     �R@      8@                      @      <@               @       @              Z@              D@      "@              "@     �P@     @c@      @      4@     �`@     �C@     @n@      I@      l@     �Z@      (@      "@     �C@      W@      @      2@      Y@      7@     �U@     �D@     �T@     @P@       @              <@      O@      �?       @      A@      0@     �c@      "@     �a@     �D@      @      0@      i@     �p@      1@      ?@     �l@     �L@     �r@      `@     �q@     �e@      5@      �?     �F@      O@       @      @      J@       @      ^@      3@      X@      <@      @      �?      D@      N@       @      @      C@       @     �[@      (@     @V@      8@      @      �?      .@      *@               @      6@       @      :@      @      3@      @      @              9@     �G@       @      �?      0@             @U@       @     �Q@      2@      �?              @       @              @      ,@              "@      @      @      @                              �?              �?      "@              "@      @      @       @                      @      �?               @      @                       @      �?       @              .@     `c@     �i@      .@      9@     @f@     �K@     @f@     �[@     �g@      b@      1@       @     �a@      h@      ,@      9@     �d@     �H@      f@     �X@      f@     ``@      ,@      @      Z@     @`@      $@      0@     �[@      E@     @R@      T@      T@     �X@      *@      �?      C@     �O@      @      "@     �K@      @     �Y@      2@     @X@     �@@      �?      @      *@      (@      �?              *@      @       @      (@      &@      *@      @              @      @                      "@      @       @      @      �?      @      @      @      @      @      �?              @                      @      $@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�*�rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���D�`@�	           ��@       	                     @'���+@�            �@                           �?*�̺�@_           ��@                           �?{�&ѧ>@*            }@������������������������       ����֐@F            �\@������������������������       �m��.Mg @�            �u@                           @H_��Ҫ@5           ��@������������������������       �Ls��@A           `}@������������������������       ���YE�T@�             x@
                           �?���GS@8           `}@                           @���@�            @o@������������������������       �Of3��)@@            @Y@������������������������       ��$lѰ�@a            �b@                           @�)k$@�            �k@������������������������       �0��R(@3            �Q@������������������������       �}_�pB@d            �b@                           @� &�0�@#           ��@                          �6@�v��	@;           P�@                           �?tk9@��@�            �x@������������������������       ���5DPi@c            �b@������������������������       �S$�wd�@�             o@                          �8@�mEPv�	@=           (�@������������������������       �Ϭr���@�            �q@������������������������       �y����	@�           H�@                          �6@U'_���@�           ��@                           @N]��S@�            �r@������������������������       �L:���@&             P@������������������������       �S��[@�            `m@                           @��].�I@3           P�@������������������������       ���ɮ�@�             t@������������������������       ���r��@t             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �q@     @�@      B@      J@     �z@     @Z@     t�@     @j@     8�@     w@      >@      @     @V@     �m@      ,@      ,@      d@      7@     ȃ@      S@     �x@      a@      @      �?      P@     �e@      "@       @     @Z@      ,@      @      N@     �q@     �Y@      @              3@      N@               @      B@       @     �j@      *@     @X@      9@                      @      4@                      2@       @      >@      @      5@      (@                      ,@      D@               @      2@             �f@      @      S@      *@              �?     �F@     �\@      "@      @     @Q@      (@     �q@     �G@      g@     �S@      @      �?     �A@     @R@       @       @      J@      (@      [@     �C@     �T@     �J@      @              $@      E@      �?      @      1@             @f@       @     @Y@      9@              @      9@      P@      @      @     �K@      "@     �`@      0@     �\@     �@@       @      @      ,@     �A@       @      @     �E@      @      G@       @      M@      9@       @      @      "@      &@      �?              @      @      7@       @      ;@      (@      �?              @      8@      �?      @      B@      @      7@      @      ?@      *@      �?              &@      =@      @      �?      (@       @     @V@       @     �L@       @                      �?      0@      @      �?       @      �?      :@      @      &@       @                      $@      *@                      $@      �?     �O@      �?      G@      @              0@     �h@     �s@      6@      C@     �p@     �T@     @z@     �`@     �w@      m@      8@      0@      c@      j@      1@      A@      f@      M@      g@     �W@     @f@     `d@      4@      @     �K@     @T@      @      .@     �D@      3@     @Q@      7@     �M@      =@              @      9@      >@      @      @      (@      @      C@       @      0@      *@               @      >@     �I@              &@      =@      .@      ?@      5@     �E@      0@              &@     @X@     �_@      ,@      3@     �`@     �C@     �\@     �Q@     �]@     �`@      4@             �B@     �@@      @      $@      J@       @     �E@       @      E@      D@      @      &@      N@     �W@      "@      "@     �T@      ?@      R@     �O@     @S@     �W@      ,@              F@     @Z@      @      @      V@      8@     �m@      D@      i@     �Q@      @              "@     �E@      @              <@      *@     �Z@      �?     �Q@      5@      @                      (@                      $@      "@      3@      �?      "@       @       @              "@      ?@      @              2@      @     �U@              O@      3@       @             �A@      O@       @      @      N@      &@     @`@     �C@     @`@     �H@                      3@     �B@               @      B@      @     �X@      2@     �U@      6@                      0@      9@       @       @      8@      @      @@      5@      F@      ;@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ_��mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�׳D��@�	           ��@       	                    �?�d�*̎	@           (�@                           �?��Q�9�@6           �}@                          �7@1�q�6@�            �k@������������������������       ���՜&@Y            �`@������������������������       ���H�[1@8             V@                           �?t�.L�]@�            �o@������������������������       ��me�P@D            �W@������������������������       �ݺ�Zu@a            �c@
                           �?���n0
@�           ��@                          �?@�+��)@           y@������������������������       �@r��H�@�             x@������������������������       ���qa@	             .@                            �?�.F�i
@�           ��@������������������������       �Èe���@�            �l@������������������������       �u�Hm	�
@C           �@                          �2@�ao^��@�           ��@                           @���0�@�           ؆@                            �?Fb�l��@k            @e@������������������������       ���G@2            @T@������������������������       �vZ�7�@9            @V@                          �1@:�R�� @`           ��@������������������������       ���0V^��?�            �v@������������������������       �y�V��@�             i@                           �?����@�           ��@                           �?�'K~@'           �}@������������������������       � n�+J@�            �q@������������������������       ��#�5@w            �g@                          �7@w�b{�@�           �@������������������������       �Og?(1_@�           ؄@������������������������       �J�J5@           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@      �@     �C@     �L@     �}@     �S@     p�@     �m@     x�@     �w@     �B@      *@     �e@     @l@      ?@      D@     �o@     �G@      h@     �`@      p@     @j@      @@              F@     �R@      @      @      M@      @     �T@     �A@     �Z@      K@      @              0@      A@      @      @      <@      @     �F@      2@      E@      6@       @              $@      ,@                      3@       @     �C@      *@      9@      "@       @              @      4@      @      @      "@      �?      @      @      1@      *@                      <@      D@              �?      >@              C@      1@      P@      @@      @              $@      &@                      "@              6@      @      <@      "@       @              2@      =@              �?      5@              0@      *@      B@      7@      �?      *@      `@      c@      :@     �@@     �h@      F@     �[@      Y@     �b@     �c@      ;@      �?      :@     �Q@      @      ,@     �T@      @     �K@      >@      B@     �Q@      @      �?      7@     �Q@      �?      ,@      T@      @     �K@      ;@     �A@     @Q@      @              @              @              @                      @      �?      �?              (@     �Y@     @T@      5@      3@     �\@     �C@     �K@     �Q@     �\@     �U@      6@             �E@      2@       @      @      G@      "@      "@      @@      =@      7@      .@      (@     �M@     �O@      3@      .@      Q@      >@      G@      C@     @U@     �O@      @             @_@     �s@       @      1@     �k@      @@     h�@     �Y@     x�@      e@      @              5@     �W@       @      @      A@       @     �u@      :@      d@     �C@      �?               @      ;@              @      *@      �?      L@      0@     �B@      .@                       @      3@                      @      �?      :@      @      ,@       @                               @              @      "@              >@      "@      7@      @                      3@     �P@       @       @      5@      �?     0r@      $@     �^@      8@      �?               @     �D@               @      2@             �h@      @     �S@       @      �?              &@      :@       @              @      �?      W@      @     �F@      0@                      Z@      l@      @      (@     @g@      >@      {@      S@     �v@      `@      @              2@      P@      �?      �?      D@      @     �f@       @     �`@      9@      �?              *@     �A@              �?      <@      �?     �_@      @     �N@      0@                      @      =@      �?              (@      @      K@      @     �Q@      "@      �?             �U@      d@      @      &@     @b@      7@     �o@      Q@     `m@      Z@      @             �F@     �Z@      @      @     @U@      *@     @g@      =@      `@     �N@       @             �D@      K@      �?      @     �N@      $@     �P@     �C@     �Z@     �E@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@V@�	i@�	           ��@       	                    �?�� f�@~           :�@                           @-�1p�@�           �@                           �?i�
]�a@�            �v@������������������������       ������@�            �o@������������������������       ��R�8�@H            @\@                           �?S&R9�Z�?�            �v@������������������������       ������?�             h@������������������������       �?w.=�?n            �e@
                          �1@5�9r�@�            �@                           @x�O��)@�            0w@������������������������       �\��}� @"             I@������������������������       ����E�@�            t@                           �?�A��<]@�           4�@������������������������       ���,�i@4            �V@������������������������       ��tЎ[@|           ��@                           �?���u��@R           ��@                           �?! �[(@1           �}@                           �?J��"�	@�            `n@������������������������       �aO��+�@6            �V@������������������������       ��H��{*@f             c@                            @i�6�@�             m@������������������������       �Ŷ"�4n@v            �e@������������������������       �ANbx�)�?            �M@                           �?�&�4<�	@!           @�@                           �?k����@A            @Y@������������������������       ��eO���@'            �O@������������������������       ���"��@             C@                            �?���*�r	@�           ��@������������������������       ��C�[�	@w           8�@������������������������       ����@i            �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      s@     �@      ;@     �R@     �z@     �U@     ��@     `i@     ��@     Px@      @@       @     �_@      s@      $@      =@      i@      ;@      �@     �W@     �@      f@      &@              C@     @U@              @     �F@       @     ps@      <@     �e@      F@       @              :@      E@              @     �@@       @      [@      8@     @W@      A@      �?              1@     �@@               @      7@       @     @R@      2@     �K@      >@      �?              "@      "@               @      $@             �A@      @      C@      @                      (@     �E@              �?      (@             `i@      @      T@      $@      �?               @      3@              �?       @              \@      �?     �B@      @                      @      8@                      @             �V@      @     �E@      @      �?       @     @V@     `k@      $@      8@     �c@      9@     �x@     �P@      u@     �`@      "@      �?      2@     �N@      �?      @      :@      �?     ``@      &@     �U@      =@                      @                              �?              8@       @      @      @              �?      &@     �N@      �?      @      9@      �?     �Z@      @     @T@      9@              @     �Q@     �c@      "@      3@     @`@      8@     �p@      L@      o@     �Y@      "@       @      �?      1@              @      1@      @      @       @      5@      "@              @     �Q@     �a@      "@      ,@     @\@      4@     @p@      H@     �l@     �W@      "@      (@      f@     @j@      1@     �F@     �l@      N@      s@      [@     `s@     �j@      5@             �C@     @P@       @      @      K@      @      ]@      2@      ]@     �K@      @              <@     �E@       @      @      C@       @     �@@      @      I@     �A@       @              ,@      $@                      *@              7@              2@      (@      �?              ,@     �@@       @      @      9@       @      $@      @      @@      7@      �?              &@      6@                      0@      @     �T@      &@     �P@      4@      �?              "@      6@                      *@      @      I@      @      K@      .@      �?               @                              @             �@@      @      (@      @              (@     @a@      b@      .@      E@     �e@     �K@     �g@     �V@     @h@     �c@      2@      @      5@      @              "@      2@      @      @      1@      &@      @              @      0@      @               @      ,@      @      @      @      @      @                      @      @              @      @      �?      �?      $@      @       @               @     @]@     `a@      .@     �@@     �c@     �I@     @g@     @R@     �f@     �b@      2@      @     �R@     @P@      @      1@      Q@      =@     �W@     �H@      U@     �S@      ,@      @     �E@     �R@      $@      0@     @V@      6@     �V@      8@     �X@     @R@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJR�
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��w&�%@�	           ��@       	                     @ќi7F@c           2�@                           �?W��@�           D�@                           @��ᔞ�@l           Ȃ@������������������������       �n����@�             o@������������������������       ��R�]�?�            v@                           @���@�           ��@������������������������       �������@           `|@������������������������       �^��,��@q           ��@
                           �?^�[�Q�@i           @�@                          �1@�F�SI@�            �s@������������������������       ��`���@,            @R@������������������������       ����"ڇ@�            �n@                           @˽ T��@�            �p@������������������������       �8���:�@5            @T@������������������������       ��/&�:@q             g@                           @�.�q�@S           ��@                           �?
�cx�	@�           �@                           �?�z�+@�             r@������������������������       �;���3�@^             b@������������������������       �����Z@_            �a@                           �?��E�
@           Ȉ@������������������������       ����~`�@,             O@������������������������       �@�//��	@�           ؆@                          �6@}ِ@�           ��@                            @)+��=z@H            @\@������������������������       �} ��@8             W@������������������������       �������?             5@                           @����B@B           0�@������������������������       ���֟��@�            �t@������������������������       ��w��@x            @g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     s@     ��@     �C@     �P@     �y@     �R@     d�@     �g@     ؊@     pt@      @@      @     @^@     �s@      0@      @@      h@      5@     ��@      T@     h�@      b@      $@      @     �T@     �m@      @      5@     �`@      "@     ��@      P@     0x@     �X@      @              >@     �S@      �?      �?      =@       @     �p@      &@     �b@      =@       @              1@      7@      �?              0@      �?     �T@      @     @S@      6@       @              *@      L@              �?      *@      �?     @g@      @      R@      @              @      J@     �c@      @      4@     �Z@      @     �r@     �J@     �m@     �Q@      @      @     �@@     �R@      @      $@      Q@      @     �X@      F@     �R@     �A@      @              3@      U@              $@      C@       @     @i@      "@     `d@     �A@              @     �C@      T@      $@      &@     �L@      (@     �d@      0@     @a@     �F@      @      @      ?@      G@       @      @      E@      "@      P@       @     �O@      B@      @              "@      @      �?      �?      @              ?@       @      @      &@              @      6@     �C@      @      @     �B@      "@     �@@      @     �L@      9@      @               @      A@       @      @      .@      @     �Y@       @     �R@      "@       @              @      0@              @       @       @      ;@      @      1@      @                      @      2@       @       @      *@      �?      S@      @      M@      @       @      *@      g@      l@      7@      A@      k@      K@     �s@     �[@     �t@     �f@      6@      *@     @b@     @a@      ,@      9@     �c@     �F@      a@     @W@      d@     �`@      5@       @      @@     �D@      �?      @     �B@              P@      &@      N@      =@      @       @      2@      9@      �?      @      ,@             �A@      @      7@      2@                      ,@      0@              �?      7@              =@      @     �B@      &@      @      &@     �\@     @X@      *@      3@      ^@     �F@     @R@     �T@      Y@     �Y@      0@       @      *@      @               @      (@      �?      �?      @      "@      @      @      "@     @Y@     �V@      *@      1@      [@      F@      R@      S@     �V@     �X@      $@              C@     �U@      "@      "@     �M@      "@      f@      1@     �e@     �I@      �?              @      &@       @              $@      @     �F@              3@      &@                      @      "@       @              $@      @     �D@              @      $@                               @                                      @              ,@      �?                      @@      S@      �?      "@     �H@      @     �`@      1@     `c@      D@      �?              0@      I@              @      >@       @     @X@      @      Z@      8@      �?              0@      :@      �?      @      3@      @     �A@      (@     �I@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Ї�T�@@�	           ��@       	                    �?��j���@y           X�@                           �?2�vA	@           @�@                            �?�a��S	@|           ��@������������������������       �)H�d@�            s@������������������������       ��dz��J	@�            @t@                            �?$Իd@�            `n@������������������������       ���2R�@0            �Q@������������������������       �U��W�@l            �e@
                          �1@W��Єy@a           �@                          �0@�s���@l            @e@������������������������       �pȇ�9@!             K@������������������������       ��K
�,�@K             ]@                           �?R�(;��@�           h�@������������������������       �YƥC�@�            q@������������������������       �u�3GQ	@D           H�@                           �?&��B�@#           t�@                           �?f�S^c� @\           `�@                          �3@h�q*f[ @�             u@������������������������       ���;T���?u            @h@������������������������       �A��Rܮ @]             b@                          �8@�M��?@�            @k@������������������������       ��I��5� @w            `g@������������������������       �`�dR]��?             ?@                           @M-�`�@�           đ@                           �?r,��?}@�           L�@������������������������       �-�.ւ@R           0�@������������������������       �m?��@@a           h�@                           @ܣr�`�	@             >@������������������������       �j{��0J@             *@������������������������       ��{�V�@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pr@     �@      :@      E@     @~@     �V@      �@     @j@     ��@     �v@      :@      6@     �k@     0v@      3@      =@      u@     @S@     0v@     `e@     �v@     @n@      8@      *@     �V@      c@      *@      $@      ^@      D@      a@      Q@     @_@     �X@      @      *@     @P@      _@      (@      @     �W@      =@     �S@      H@      S@     @S@      @      @      >@     @S@      @      �?     �C@      .@      G@     �A@      9@      :@      @      $@     �A@     �G@       @      @     �K@      ,@     �@@      *@     �I@     �I@      �?              9@      <@      �?      @      :@      &@      M@      4@     �H@      6@                       @      .@              �?      "@              6@      @      $@      @                      7@      *@      �?       @      1@      &@      B@      ,@     �C@      1@              "@     �`@     `i@      @      3@     @k@     �B@     @k@     �Y@      n@     �a@      3@              @      @@              �?      7@              I@      @     �E@      $@                       @      .@              �?      $@              ,@      �?      @      @                      @      1@                      *@              B@      @     �B@      @              "@     @_@     `e@      @      2@     `h@     �B@      e@     �X@     �h@     �`@      3@              @@      F@              �?      =@      �?      L@      &@      Q@      ?@              "@     @W@     �_@      @      1@     �d@      B@      \@      V@     @`@     �Y@      3@             @R@     �k@      @      *@     @b@      ,@     �@     �C@     `z@     �]@       @              2@      S@      �?      �?      C@      �?     �p@      @      _@      6@                      &@      E@              �?      :@             �e@       @     �Q@      ,@                      "@      1@              �?      &@              Y@             �I@      @                       @      9@                      .@              R@       @      3@      "@                      @      A@      �?              (@      �?     �X@      @      K@       @                      @      @@      �?              "@             �W@      @     �A@      @                               @                      @      �?      @              3@       @                     �K@     @b@      @      (@      [@      *@     �v@      A@     �r@      X@       @              J@     �a@      @      "@      Z@      $@     �v@      @@     pr@     @W@       @              ;@      T@       @       @      N@       @     @c@      &@     �`@     �G@      �?              9@      O@      @      @      F@       @      j@      5@     `d@      G@      �?              @      @      �?      @      @      @      @       @      @      @                      �?              �?              @       @               @      �?      @                       @      @              @      �?      �?      @               @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ"�K hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ݨ�
�g@�	           ��@       	                    @�"���@           ��@                          �;@Ix��B(@�           ��@                           �?�l��@y           ��@������������������������       �5����X@�            @r@������������������������       ��U�' @�            s@                            �?$�V�@7            @X@������������������������       �4�-Z�@            �E@������������������������       ��Iۜt@             K@
                          �4@9�&#^ @a           Ё@                           @{���
3�?�            �w@������������������������       �͌����?�            �k@������������������������       ���w#1 @c             d@                          �8@�u5��@~            �g@������������������������       �`����@Q             _@������������������������       �k�m�T@-             P@                            �?N�1�w@�           ��@                           �?��:�f�@�            �@                           �?�YtH�	@�            �t@������������������������       �ġj�@S             _@������������������������       ������2	@�            `j@                          �6@�o��lo@�            Pu@������������������������       �Йx	��@�            �i@������������������������       �4�w��;@X             a@                           @I5�j�U@�           Ԟ@                          �?@e��D~	@�           �@������������������������       �I�4`	@�           p�@������������������������       �m���8@            �D@                          �<@t����@4           ��@������������������������       ��׏,o1@           ؉@������������������������       ��^_׍�@#            �J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �s@     8�@      ;@      M@     �{@      U@     �@     �k@     ��@     �w@     �A@      @     �R@     `d@      �?      *@      ]@      @     @      F@     �p@     @T@      @      @     �L@     �V@      �?      *@      U@       @     `i@      B@      b@     �L@      @              D@     �T@      �?      @     �Q@       @     @h@      9@     ``@      E@       @              .@      B@      �?      @     �D@       @     @Z@      2@      I@      0@      �?              9@     �G@                      =@             @V@      @     @T@      :@      �?      @      1@       @              @      ,@              "@      &@      *@      .@      �?      @      @      �?              @      @              �?      @      @      ,@      �?              &@      @              @      $@               @      @       @      �?                      1@      R@                      @@      @     `r@       @      ^@      8@                      *@      B@                      0@             �k@      @     �S@      *@                       @      8@                       @              a@      �?      G@      @                      @      (@                      ,@             @U@       @     �@@      $@                      @      B@                      0@      @      R@      @     �D@      &@                      @      <@                      (@             �G@              ;@      @                               @                      @      @      9@      @      ,@      @              1@     �m@     @v@      :@     �F@     pt@     �S@     ��@     `f@     X�@     �r@      @@      �?     �Q@      W@      @      1@     �V@      5@     �a@      K@     �Z@      Q@      "@      �?     �F@      C@      @      *@     �O@      0@      ?@     �F@      A@     �B@       @              "@      &@              "@      6@      @      6@      ,@      3@      *@       @      �?      B@      ;@      @      @     �D@      *@      "@      ?@      .@      8@      @              9@      K@       @      @      <@      @     �[@      "@      R@      ?@      �?              "@      9@       @      �?      1@             @U@      @     �G@      *@                      0@      =@              @      &@      @      9@      @      9@      2@      �?      0@      e@     �p@      4@      <@     �m@      M@     0x@     @_@     z@     �l@      7@      0@     @]@     �c@      *@      1@     �a@     �G@     �`@     @Z@      f@     @c@      .@      (@      Z@     �b@      &@      1@     `a@     �F@     �`@     @Z@     �e@      b@      .@      @      *@      @       @              @       @                       @      "@                      J@     �Z@      @      &@     �W@      &@     �o@      4@      n@      S@       @             �E@     �Z@      @      $@      S@      &@     �n@      4@     `m@     @P@       @              "@      �?      �?      �?      2@              @              @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>�0\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����Q@�	           ��@       	                     �??Q�Y��	@�           8�@                          �:@�����D	@>           �@                           �?r���y�@            y@������������������������       ��Ԅ���@j            �e@������������������������       ��
pɭ@�            �l@                           �?v�� 	@;            �Y@������������������������       �Bmֺ�@             :@������������������������       ����z3	@+             S@
                           �?��/,7�	@�           X�@                           @hkx)�	@           �x@������������������������       �
��O�	@�            �v@������������������������       �T�\>�@             9@                           �?�q��	@�           p�@������������������������       ���y���@�            @o@������������������������       �DoR_
@%           @}@                          �5@��Ԝz@�           ��@                           �?e��c��@�           4�@                          �3@'|�` @V           H�@������������������������       ��m"��?�            px@������������������������       �q>_$= @_            @d@                          �4@0E����@5            �@������������������������       ���}�"�@�           x�@������������������������       �] z-b�@Z            �b@                           �?��j��@           p�@                           @T{1y�7@�            �k@������������������������       ����5�@Q            �_@������������������������       �Jn��@?             X@                           @|F��f=@�           x�@������������������������       ����'�@u             e@������������������������       ��y��f@           `z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     0r@     ؀@     �@@     �K@      {@     �T@     ��@      n@     �@     �v@      8@      :@      e@     `l@      <@      D@     @m@     �H@     �l@     �b@     �m@     �i@      4@      @      L@     �S@      @      3@     �Q@      &@      R@      H@     �T@     �I@      @      �?     �I@      Q@      @      0@     �M@      @     �O@     �B@      P@      =@      @              $@      2@               @      <@      @     �D@      2@     �A@      &@              �?     �D@      I@      @       @      ?@      @      6@      3@      =@      2@      @      @      @      &@      �?      @      &@      @      "@      &@      2@      6@       @      @              @                      @      �?      @      @       @      �?              �?      @       @      �?      @       @      @      @       @      $@      5@       @      5@     @\@     �b@      7@      5@     �d@      C@     �c@     @Y@     @c@     `c@      ,@       @     �G@     �M@      (@       @      J@      *@     �K@      @@     �G@      L@      @       @     �G@     �J@      (@       @     �F@      &@     �K@      ;@     �G@     �I@      @                      @                      @       @              @              @              *@     �P@     @V@      &@      *@      \@      9@     �Y@     @Q@     �Z@     �X@      &@      @      4@     �B@               @      F@      �?      J@      1@     �F@      <@      �?      $@      G@      J@      &@      &@      Q@      8@     �I@      J@      O@     �Q@      $@      �?     �^@     �s@      @      .@     �h@     �@@     �@     �V@     ��@     @c@      @              M@     �j@       @      @     �W@      (@     @�@     �A@     �v@      U@      @              7@     �O@              �?      <@              r@      @      _@      3@       @              2@      C@                       @             �i@      @      Y@      1@       @              @      9@              �?      4@              U@      �?      8@       @                     �A@     �b@       @      @     �P@      (@     �t@      >@     �m@     @P@       @              >@      ^@       @      @     �J@      @     �r@      <@     @g@     �K@                      @      =@              �?      ,@      @      >@       @      I@      $@       @      �?      P@      Y@      @       @     �Y@      5@     `k@      L@      e@     �Q@                      "@      >@      �?              2@      @     �S@      $@      L@      ,@                      "@      0@                      @      @      I@      @      A@       @                              ,@      �?              (@              =@      @      6@      (@              �?     �K@     �Q@       @       @     @U@      .@     �a@      G@     @\@      L@                      6@      8@              @      ;@      @      8@      5@      3@      6@              �?     �@@      G@       @      @      M@       @      ]@      9@     �W@      A@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B                             �?�2���@�	           ��@       	                    �?���Z@'           `�@                            @/���@5           ~@                           �?.z�@�            �p@������������������������       �o��͝�@X            @a@������������������������       �F���I�@^             `@                           �?��Œ@            �j@������������������������       ��c���{@>            @[@������������������������       �e�rIq@A            �Z@
                          �=@d��X@�           ��@                           �?�[��}�@�           @�@������������������������       �^b8��@            {@������������������������       �Y=	��@�            `s@������������������������       �1�����@             .@                           !@�E-�j@�           �@                           @x��K�X@�           ��@                           �?�2O]�	@�           ��@������������������������       ����]B
@�           đ@������������������������       �.�c��K@           @{@                          �4@L��sȏ@�           ̐@������������������������       ��&I(@X           ��@������������������������       �=��g�A@V           ��@������������������������       ��B�:��@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     X�@      ;@     @R@     �{@      V@     x�@     @l@     Ј@     �u@      F@      �?      T@     �e@      @      1@     @[@      &@     `z@     �B@     �q@     @W@      @      �?     �G@     �T@       @      ,@     �N@      @     @W@      <@     �W@     �I@      @      �?      =@      @@      �?      @     �B@      �?      M@      "@      M@      @@      @      �?      .@      *@                      6@              A@      @      @@      0@      �?              ,@      3@      �?      @      .@      �?      8@      @      :@      0@      @              2@      I@      �?      $@      8@      @     �A@      3@      B@      3@                      @      5@      �?      @      0@      @      6@      @      5@      @                      &@      =@              @       @              *@      *@      .@      ,@                     �@@     �V@       @      @      H@      @     �t@      "@      h@      E@      @              @@     �V@       @      @     �F@      @     `t@      @     �g@      E@                      (@     �J@              @     �A@      @      i@      @      X@      =@                      4@     �B@       @              $@      @     �_@      @     �W@      *@                      �?                              @      �?      @       @       @              @      4@     �i@     �w@      7@      L@     �t@     @S@     H�@     �g@     �@     p@     �B@      4@     @i@     �w@      7@      L@     `t@     �R@     H�@     �g@     �@     �o@      @@      3@     �a@     �k@      1@      F@     �l@      P@      l@     �e@      m@     `f@      :@      3@      Z@     `c@      1@      C@      e@     �K@     @a@     �`@      c@     �`@      9@              B@      Q@              @      O@      "@     �U@     �D@      T@      G@      �?      �?      O@     �c@      @      (@      X@      $@     �v@      .@     q@      S@      @              :@     @R@       @      @      =@      �?     �l@      @      a@     �B@              �?      B@     @U@      @      @     �P@      "@     �`@      (@      a@     �C@      @              @       @                       @      @                       @       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��+"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����1@�	           ��@       	                    �?�RE���@�           >�@                          �;@��LP�	@           h�@                           �?aR��@f           `�@������������������������       ��� �"�@           pz@������������������������       ��+���Q	@[           ��@                           �?g����	@�             p@������������������������       ���` @#            �K@������������������������       �N|r��x	@�            `i@
                          �4@`��@z           (�@                           �?��vy)D@�            �r@������������������������       ��(4��@J            �\@������������������������       ��~��A@p            �f@                           �?�Ki
s�@�            �q@������������������������       �jG'|b�@2             U@������������������������       �(��|.@�             i@                          �4@8�	��@>           ��@                           @0��З@G           0�@                          �1@�Wl��@�             i@������������������������       �fu��_��?4            �T@������������������������       �tIi�N|@M            �]@                            �?H���� @�           ��@������������������������       ��;����?b             b@������������������������       �����>l@d           h�@                           @#�y}�@�            �@                            @U�.�i@E           �@������������������������       �3�y��@           �{@������������������������       ��p �f�?(            �Q@                          �7@��XNG@�            0r@������������������������       �{e��MJ@M            @_@������������������������       �"p	�D@e            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     `r@     ��@     �@@     �F@     �|@     @R@      �@     �j@     ��@     @w@     �B@      (@     @j@     �t@      5@     �B@     Pt@      L@     �x@     @f@     pu@     �p@      =@      (@     �d@     @o@      4@      ?@     �n@      D@     �n@      a@     `m@     �j@      <@      @      a@      l@      (@      6@     `k@      <@     �k@      \@     �j@     `b@      :@             �D@     @S@               @      I@      �?      X@      8@     @W@      B@      @      @     �W@     `b@      (@      4@      e@      ;@     �_@      V@      ^@     �[@      7@      @      =@      :@       @      "@      <@      (@      8@      9@      6@     �P@       @      �?      @       @              @      @      �?      &@      @      @      (@              @      8@      2@       @      @      6@      &@      *@      6@      2@     �K@       @             �F@     @U@      �?      @     �S@      0@      b@     �D@      [@     �K@      �?              *@     �E@      �?       @      >@      @     @X@      7@      O@      6@                      @      2@      �?              2@      @      ?@       @      6@      @                      @      9@               @      (@      �?     �P@      .@      D@      .@                      @@      E@              @      H@      (@      H@      2@      G@     �@@      �?              "@       @                      *@      @      8@              4@      @                      7@      A@              @     �A@       @      8@      2@      :@      ;@      �?      �?      U@      n@      (@       @      a@      1@      �@      A@     pz@     �Y@       @             �D@      \@      @      @     �H@      @     `z@      (@     �j@     �C@                      1@      @@                      @      @      U@      @      E@       @                      @      &@                       @              F@              2@      @                      *@      5@                      @      @      D@      @      8@      @                      8@      T@      @      @     �E@              u@      @     �e@      ?@                      @      $@                      *@             �V@              6@      @                      4@     �Q@      @      @      >@              o@      @     �b@      9@              �?     �E@      `@      @      @     �U@      (@     @k@      6@      j@      P@       @      �?      7@     @S@      �?             �K@      @     �d@       @     �`@     �@@       @      �?      4@     @S@      �?              I@      @     �`@       @     �[@      ?@      @              @                              @              ?@              9@       @      @              4@     �I@      @      @      @@      @     �J@      ,@     �R@      ?@                      @     �B@      �?      @      *@      @      9@       @      ;@      $@                      0@      ,@      @       @      3@       @      <@      (@     �G@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@g�=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�ߌ�@�	           ��@       	                    �?�B�/�@2           ��@                          �<@a�І0i@�           �@                           @����}�@           ��@������������������������       � 1�HH�@�            Pu@������������������������       ��'>�2�?�            �o@                          �>@���[@            �D@������������������������       �T�48D@             7@������������������������       �2����@             2@
                          �3@��u9�@�           ��@                           @���NΎ@�            px@������������������������       �.���E@�             i@������������������������       �)�@ @o            �g@                            �?."�m��@�           �@������������������������       �\�}�N�@�            �u@������������������������       �#���#�@�            pt@                            @���׿M@�           D�@                           �?/�~U@�           ��@                           �?�wz�@           �y@������������������������       ���Ց��@e            `d@������������������������       �$�7a�(@�             o@                          �9@�Ճ���@�           ��@������������������������       ��L[�@F           ��@������������������������       �'���L�@�            �l@                           @sq�"x�@�            �@                          �7@�x���O@D           �@������������������������       �Tq�5�@�            Pu@������������������������       ��_	��@m            @e@                          �7@���c�@d            �d@������������������������       �6��^���?C            @\@������������������������       �T��@qt@!             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@     p�@      7@      M@     �{@     @S@     D�@     `m@     @�@     �v@      6@      @      ^@     �o@      @      =@     `h@     �A@     �~@      S@     �t@      c@      $@              I@     @U@      �?      (@      H@       @     �o@      8@     @^@     �A@                      H@     �S@      �?      "@      G@       @      o@      3@      \@      :@                      <@      K@      �?      @      C@       @     �Y@      .@     �P@      6@                      4@      8@              @       @             @b@      @     �F@      @                       @      @              @       @              @      @      "@      "@                              @              �?      �?              @              @      @                       @                       @      �?              �?      @      @      @              @     �Q@      e@      @      1@     `b@      ;@     �m@      J@      j@     �]@      $@      �?      6@     �J@              �?      B@      @     @a@      1@     �U@     �@@      �?      �?      (@      B@                      9@      @     �K@      ,@      <@      9@      �?              $@      1@              �?      &@             �T@      @      M@       @              @      H@      ]@      @      0@     �[@      8@     �X@     �A@     �^@     @U@      "@              ?@      P@              @     �H@      (@     �I@      :@      Q@      B@      @      @      1@      J@      @      (@      O@      (@     �G@      "@      K@     �H@       @      "@     @f@      q@      1@      =@     @o@      E@     @�@     �c@     �}@     `j@      (@      @     @[@     @f@      .@      2@     �d@     �@@      y@     �Y@     �u@     �b@      @              =@     �I@              �?      @@      @     @_@      $@     @`@      =@       @              8@      5@              �?      3@             �@@      @      H@      *@      �?              @      >@                      *@      @      W@      @     �T@      0@      �?      @      T@     �_@      .@      1@     �`@      >@     Pq@      W@     �k@      ^@      @      @      L@     �[@      *@      *@      X@      2@     0p@     �L@     �f@     �T@      @       @      8@      1@       @      @      C@      (@      2@     �A@      C@      C@              @     @Q@     �W@       @      &@      U@      "@     �b@     �L@      `@      O@      @      @      J@     �U@      �?      $@     @R@      @     �T@      L@     @T@     �J@      @      @      ;@      M@              @     �E@       @      J@      @@      R@      E@      @              9@      <@      �?      @      >@      @      ?@      8@      "@      &@       @              1@       @      �?      �?      &@      @     �P@      �?     �G@      "@                      "@      @                      @      @      K@              A@      @                       @      @      �?      �?       @              *@      �?      *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ\��VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�w��@	           ��@       	                   �3@�T�V�@<           �@                            �?�y;
w�@�           ��@                           �?/��'��@�            �k@������������������������       ��s�^�@4             U@������������������������       �OY'W�D@T            `a@                           �?�m�R9@1           �@������������������������       �P��E�-@\            �b@������������������������       �Z�n�@�            0v@
                           �?�w�	�/	@�           ��@                          �<@𿠊�G@�            �x@������������������������       �n���@�            @u@������������������������       ��9n�o@&             L@                           @-�U|��	@�           ��@������������������������       �5<���	@<            �@������������������������       �xͦ'	@Y            �@                           �?��[�@C           �@                            �?<6S�� @d           ��@                           �?>9���?S            �^@������������������������       �y(�[�P�?(             L@������������������������       �f�[�-� @+            �P@                          �5@R���� @           �{@������������������������       �`;{�=�?�            �r@������������������������       ���9v�@S            �a@                           @;��J�?@�           @�@                          �1@��1@           X�@������������������������       ��u4z�?a            `d@������������������������       ����1�	@�           @�@                          �5@�<��3@�            Pt@������������������������       �^�]�d�@q            �f@������������������������       ���	���@[             b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     Ps@     ��@      =@      L@     �z@     �S@     T�@     @j@     P�@     �u@      :@      $@     �j@     �u@      5@     �F@     `r@      N@     0x@     �e@     �x@      j@      7@      �?      C@     �Y@      @      &@     �V@      (@     �f@      G@     �e@      P@      @              @     �C@                      2@      �?     �M@      (@     �Q@      ,@       @                      3@                      @              ;@       @      6@      �?                      @      4@                      &@      �?      @@      @     �H@      *@       @      �?      ?@     �O@      @      &@      R@      &@      _@      A@     �Y@      I@      �?              $@      9@                      0@             �F@      *@      <@      &@      �?      �?      5@      C@      @      &@      L@      &@     �S@      5@     �R@     �C@              "@     �e@     �n@      2@      A@     �i@      H@     �i@     �_@      l@      b@      4@             �F@     @R@       @      @      F@      @     �Y@      4@     �R@      9@       @             �D@     @P@       @              @@      @     �X@      .@     @Q@      *@      �?              @       @              @      (@              @      @      @      (@      �?      "@      `@     �e@      0@      >@      d@     �F@     @Y@     �Z@     �b@     �]@      2@      "@     �J@     �Q@       @      *@     �V@      ;@     �L@     �C@     �P@      R@      @              S@     �Y@       @      1@     �Q@      2@      F@     �P@     �T@     �G@      (@             @X@     �n@       @      &@     �`@      3@     ��@      C@     �w@     �a@      @              ,@     @U@      �?              >@       @     �q@       @     �[@      @@      �?                      0@      �?               @       @     �P@              4@      $@                              @                       @      �?      @@              *@      @                              (@      �?              @      �?      A@              @      @                      ,@     @Q@                      6@              k@       @     �V@      6@      �?              &@     �I@                      ,@             �d@      @     �H@      @      �?              @      2@                       @             �I@       @      E@      1@                     �T@      d@      @      &@     @Z@      1@     �w@      >@     �p@      [@       @              H@     �[@       @      @     @Q@      (@     s@      3@     �i@      O@       @                      ,@                      "@             @T@              G@      *@                      H@     @X@       @      @      N@      (@      l@      3@      d@     �H@       @             �A@     �H@      @      @      B@      @     �Q@      &@      O@      G@                      .@      ;@       @      �?      5@              O@      @      <@      5@                      4@      6@      @      @      .@      @      "@      @      A@      9@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ7�}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@'��" y@�	           ��@       	                    �?f୦��@�           4�@                            �?	{���@.           p}@                          �2@L$���3@T            �`@������������������������       ��0=�g@8            �U@������������������������       �e�1U/�@            �G@                          �2@w\��J@�             u@������������������������       �
����@�            @j@������������������������       �U��_t?	@K             `@
                           @�XЃ	@k           ��@                           @@<�\cj@�           `�@������������������������       �`0��p@�            �q@������������������������       �T/F�ڵ @�            �x@                           @68Oa=�@�            �t@������������������������       �h^vg��@L            �`@������������������������       �k����@u            �h@                           �?�j���@           ��@                           �?��6���	@�           4�@                          �9@��� �@	           @y@������������������������       �)(�0�[@�            @r@������������������������       ��cG�D	@N             \@                           �?j�Q7��	@�           ȇ@������������������������       ���:�	S
@�            q@������������������������       �� 5Q}L	@-           �~@                          �<@P���@7           ��@                           @���0p'@�           ԑ@������������������������       �	ٵ�O�@�           ��@������������������������       ����j��@N            �_@                            �?�U��p@J            �^@������������������������       �	�!Wj@             =@������������������������       ����V@6            @W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     Ȁ@      :@      P@     P@      U@     X�@      k@     ��@     �v@      A@      @     @Q@     �h@      �?      0@     @`@      ,@      �@     �O@     pt@     �]@      �?      @      <@      N@      �?      &@     �S@      *@     �Y@      >@      T@      O@      �?               @      3@                      7@       @      ?@      (@      >@      ,@                       @      2@                      *@       @      5@      @      5@       @                              �?                      $@              $@      @      "@      (@              @      :@     �D@      �?      &@      L@      &@     �Q@      2@      I@      H@      �?      �?      2@      ;@              @      F@      �?     �F@      $@     �@@      8@              @       @      ,@      �?      @      (@      $@      :@       @      1@      8@      �?             �D@      a@              @     �I@      �?     �{@     �@@     �n@     �L@                     �A@     �X@               @      >@      �?     �s@      3@     �c@      9@                      4@     �I@                      $@      �?     @^@      @     �O@      .@                      .@     �G@               @      4@             �h@      *@     �W@      $@                      @     �C@              @      5@             @_@      ,@     �V@      @@                      @      6@                      @             �J@      (@      ;@      "@                       @      1@              @      ,@              R@       @     �O@      7@              0@     �l@     @u@      9@      H@     0w@     �Q@     �z@      c@     �}@     �n@     �@@      .@      b@     �e@      1@     �A@      j@     �F@     @X@      W@      f@     �a@      7@       @      A@     �P@      @      (@     @Q@      &@      K@      6@     �S@     �F@      @              6@     �H@      @      &@      K@      @     �G@      *@     �P@      4@       @       @      (@      2@      �?      �?      .@      @      @      "@      &@      9@      @      *@     �[@     @Z@      *@      7@     `a@      A@     �E@     �Q@     �X@     �W@      1@      @      C@      F@      $@      &@      D@      1@      0@      7@      >@      B@      @       @     @R@     �N@      @      (@     �X@      1@      ;@     �G@      Q@     �M@      ,@      �?     �T@      e@       @      *@     `d@      9@     �t@     �N@     �r@     @Z@      $@      �?      P@     �c@      @      *@     �a@      7@     �s@     �J@     �q@     �S@       @      �?     �L@     �`@      @      (@      _@      4@     �q@     �D@     �p@     �R@      �?              @      8@      @      �?      0@      @      @@      (@      1@      @      @              3@      "@       @              7@       @      0@       @      .@      :@       @              @      @                      @      �?               @      @      @       @              .@      @       @              4@      �?      0@      @      $@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?}
T��r@�	           ��@       	                     �?�x'��@           P�@                           @Ti.�x�@�            Pu@                           �?> �/j�@            @j@������������������������       ��3�ϖB@Y            �b@������������������������       �\��ڤ@&            �M@                          �5@�гk# @Q            ``@������������������������       �E�-�<�?8            �W@������������������������       �!GW?��@            �B@
                           �?�r��{�@7           ��@                           �?[^���c@�            �w@������������������������       ���`�'�@Z             e@������������������������       �:�m��@�            `j@                            @i��on@Y            �@������������������������       ��D�E@           x@������������������������       ���'Y�N�?X            ``@                           @�!�%[@�           �@                          �4@�AԮ2�	@�           ��@                           �?l��9�@�           ��@������������������������       �����l	@            �A@������������������������       �Y�T��@p           ��@                           @*��`{
@T           ��@������������������������       �2ܽD;�	@           X�@������������������������       � �vُ�	@N            `a@                          �7@�����@�           �@                           @��/@@           �@������������������������       ���X�@           x�@������������������������       �8�FikN@
             2@                            �?RyP��@�            `p@������������������������       �z�}�N@'            �N@������������������������       �h�WFp@~             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Ps@     8�@     �C@     �E@     |@      X@     �@     �i@     8�@      w@      @@      �?     �W@     @h@      @      @     @[@      "@     py@      C@     `r@     �R@      @      �?      6@      P@      �?              A@      @     �Z@       @     @S@      3@      @      �?      6@     �I@                      7@      �?     �B@      @      I@      .@      @      �?      0@     �D@                      4@      �?      :@      @      :@      &@      @              @      $@                      @              &@              8@      @      �?                      *@      �?              &@      @     �Q@       @      ;@      @                              $@                       @              L@              7@      @                              @      �?              "@      @      ,@       @      @      �?                      R@     @`@       @      @     �R@      @     �r@      >@      k@      L@       @              F@     �M@       @      @     �H@       @     �U@      1@     �U@      <@       @              ,@      3@                      4@              J@      @      G@      (@                      >@      D@       @      @      =@       @      A@      (@      D@      0@       @              <@     �Q@               @      :@      @     �j@      *@     ``@      <@                      6@      P@              �?      6@      @     �a@      *@     �W@      6@                      @      @              �?      @             �Q@              B@      @              2@     �j@     Px@      B@     �B@     @u@     �U@     `�@     �d@     �@     Pr@      :@      2@     �b@     �m@      <@      <@     �m@     �R@      i@     �a@     �n@     �h@      9@       @      D@      T@      $@      @      X@      (@     �^@      I@      Z@      R@      @                       @              @      (@               @      @      �?      $@               @      D@     �S@      $@       @      U@      (@      ^@      G@     �Y@      O@      @      0@     �[@     �c@      2@      6@     �a@     �O@     �S@     �V@     �a@     �_@      3@      $@     �W@     �`@      0@      3@     �^@      I@      Q@      P@     @a@     �[@      0@      @      .@      6@       @      @      3@      *@      $@      ;@      @      0@      @             @P@      c@       @      "@     �Y@      (@     @v@      :@     �p@     �W@      �?              E@     �`@      @      @      Q@      $@      s@      $@      h@     �N@      �?              E@     �`@      @      @     �P@      @     �r@      $@     �g@      L@      �?                               @       @       @      @      @              �?      @                      7@      5@       @       @     �A@       @      J@      0@      S@     �@@                      @       @                      @      �?      1@      @      3@      @                      4@      *@       @       @      @@      �?     �A@      &@     �L@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�q�fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��%�a@�	           ��@       	                     �?�HB�0�@           ܓ@                           �?g3�7�@�            �t@                           �?�2���@U            �b@������������������������       �2<�[n@(             R@������������������������       ��a���i@-            �S@                          �3@X����@r            �f@������������������������       �V�Ҳ5��?>             W@������������������������       ���T��@4             V@
                           @u=�xT�@?           h�@                          �<@F��y�@#           �}@������������������������       �X�ֵ��@�            �y@������������������������       �DI)�@$            �M@                          �4@s�@           P}@������������������������       �R�_�s) @�            Pr@������������������������       �P����@m             f@                          �4@5m��VL@�           ��@                           @� �qo@�           đ@                            @��YyB%@~           �@������������������������       ��e�(G'@�            �v@������������������������       �5{���@�            �j@                           @�J5gn@j           ��@������������������������       �Ǻ"�y]@T             `@������������������������       �P��@           0{@                          �5@�)T��-	@�           ��@                           �?�y@K)�@�             o@������������������������       �b:AahZ@@            @Z@������������������������       ��~�p>@^             b@                          �9@�i���6	@!           ��@������������������������       �uIS��n@�           `�@������������������������       �E'mS�	@X           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     `s@     ��@      ;@      L@     �}@      V@     @�@     �m@     ��@      t@      ;@      @     �V@     �e@      �?      (@     @]@      &@     `|@      C@     �q@     �S@      @      @      1@      F@              @      :@      @     ``@      @     �R@      6@              @      0@      7@               @      @             �E@      @     �C@      (@              @      @      "@               @      @              9@      @      0@      @                      &@      ,@                       @              2@      �?      7@      "@                      �?      5@               @      3@      @      V@             �A@      $@                      �?      *@                      @             �F@              7@      @                               @               @      (@      @     �E@              (@      @                     �R@     @`@      �?       @     �V@      @     0t@     �@@     �j@      L@      @             �K@      P@      �?      @     �K@      @     �]@      8@     �W@      G@      @              G@     �K@      �?      @      G@      @     �]@      1@     �V@      =@      @              "@      "@               @      "@              �?      @      @      1@                      3@     �P@              �?      B@      @     �i@      "@     @]@      $@      @              ,@     �B@              �?      1@             �b@       @     �P@      @      @              @      =@                      3@      @     �K@      @      I@      @              3@     `k@     �x@      :@      F@     @v@     @S@     �@     �h@     0@     @n@      5@      @     �S@     �e@      @      *@     �\@      .@     �t@     �P@     @l@     @Z@      @      @     �J@     �V@      @      @     �T@      $@     @Z@      L@      U@     �R@      @             �A@     �J@       @              J@       @     @R@     �C@     �L@      F@      @      @      2@      C@      �?      @      >@       @      @@      1@      ;@      ?@      �?              9@      U@       @       @      @@      @     @l@      $@     �a@      >@                      (@      <@                      @      @      G@      @      :@       @                      *@      L@       @       @      =@       @     �f@      @      ]@      6@              .@     �a@     `k@      5@      ?@     @n@      O@     �j@     �`@     q@      a@      0@      @      *@     �E@      �?       @      B@      6@      >@       @     @Q@      1@      @      @      (@      =@      �?      �?      2@       @      @      @      1@      "@                      �?      ,@              �?      2@      ,@      ;@      @      J@       @      @      &@      `@      f@      4@      =@     �i@      D@      g@     @_@     �i@      ^@      (@      @     @S@     �Y@      &@      (@     �^@      ,@     �^@     �P@      ^@      N@      @      @     �I@     @R@      "@      1@     �T@      :@     �O@     �M@      U@      N@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ,�vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���?P@�	           ��@       	                    �?������@f           �@                          �0@Ils5@           Ј@                           �?%��n�@?            �V@������������������������       �7�nt @             <@������������������������       ��l���?.            �O@                            �?[���@�           ��@������������������������       �[kz�{]�?h            �c@������������������������       ��L�8��@Z           �@
                            @�����@e           ��@                           @}JF+�|@�           ��@������������������������       �4�h@           �{@������������������������       ����Q�_@h           ��@                          �3@����KU@�             w@������������������������       �H�<�A�@�            `n@������������������������       ���VAn�@N            @_@                           @�1���@L            �@                          �9@.Y�MK	@�           ,�@                           �?�k���]@|           p�@������������������������       ��m�� @            �i@������������������������       ����:@�             z@                           �?0��T��	@]           �@������������������������       �1�*�0

@           �{@������������������������       �8��I�@?            �W@                          �8@�;E��@s           �@                            �?��^q�z@�            �r@������������������������       �� �)7#@3            �S@������������������������       �2�r�Q�@�            �k@                          �:@_�CU�@�             q@������������������������       �z��1#@C            �X@������������������������       �vc��I�@m            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@      ;@      H@     ~@      W@     `�@     �h@     ��@     �u@      ?@      @     �`@     �r@      $@      2@     �k@     �C@     �@     �V@     @�@     `c@      *@              E@     @Y@      �?      @     �N@      @     �t@      6@     �g@     �B@      @                      .@                      0@             �@@      �?      4@      @                               @                      (@              @      �?       @      �?                              *@                      @              =@              (@      @                      E@     �U@      �?      @     �F@      @     �r@      5@      e@      ?@      @              �?      2@               @      @              S@      �?     �H@      @                     �D@      Q@      �?      @     �C@      @     �k@      4@      ^@      :@      @      @     �V@     �h@      "@      (@     @d@      B@     �u@     @Q@     �t@     �]@      $@      �?     �Q@      b@      @      $@     @Y@      9@     �p@     �H@     �n@     �V@      @      �?     �A@     �P@      @      @      N@      $@     �U@      A@      S@     �N@      @             �A@     �S@      �?      @     �D@      .@     �f@      .@      e@      >@      �?      @      4@      J@      @       @     �N@      &@     @S@      4@     �U@      ;@      @       @      0@     �D@               @      >@      @      M@      "@      K@      6@      @      �?      @      &@      @              ?@      @      3@      &@     �@@      @      �?      ,@     @g@     pp@      1@      >@      p@     �J@     �p@     �Z@     �t@      h@      2@      *@     �a@     �f@      (@      ;@      h@      G@     �]@     �V@      g@     �a@      .@      @     @V@      Y@      @      .@     �[@      $@     �Q@     �F@     �[@     �L@       @      @      ?@      8@      �?       @      :@              =@      @      M@      .@       @              M@      S@      @      @      U@      $@     �D@      C@     �J@      E@      @      $@     �J@     @T@       @      (@     �T@      B@     �H@     �F@     �R@     �T@      @      $@     �F@      O@       @      &@     �Q@      =@      D@      C@      J@     �R@      @               @      3@              �?      (@      @      "@      @      6@       @      �?      �?      F@     �T@      @      @     @P@      @     @b@      1@     �b@      J@      @      �?      2@      H@      @             �C@      @     �W@      @     �O@      5@      @              $@      &@      @              "@       @      :@       @       @      @              �?       @     �B@      �?              >@      @      Q@      @     �K@      ,@      @              :@      A@      �?      @      :@       @      J@      (@     @U@      ?@                       @      @      �?       @      @       @      1@      @     �G@      (@                      8@      <@              �?      3@             �A@      "@      C@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�B hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�� �H@�	           ��@       	                   �1@��J0�@h           �@                           �?k ~)(�@�           ȃ@                           �?C@�� @�            �o@������������������������       �g�᣺�@1             T@������������������������       �e��1�?p            �e@                           �?��n�@�            �w@������������������������       �bH�ہ@f             h@������������������������       �^/�kD@{            �g@
                            �?�w�@�           4�@                           �? �V{a�@*           x�@������������������������       �������@�             r@������������������������       �Ҝ8�N�@t           h�@                           �?��%(H@�           ��@������������������������       �'"Z S�@�            @k@������������������������       ����mdc@&           @|@                           �?	�����@E           �@                          �<@"�qAp�@            �|@                           �?��_�>@�            pv@������������������������       �X'U�&@z            �g@������������������������       ��'u�Xv@l             e@                           �?�R��#u@:             Y@������������������������       ���nc�@#            �N@������������������������       ����^�@            �C@                           @�Qu:X	@%           ��@                           @�^tQ�	@           `�@������������������������       ���",u	@           0�@������������������������       �P`�@             C@                           @���@           �z@������������������������       ���_ٟ�@           �y@������������������������       ��3����?
             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �s@     Ѐ@      8@     �P@     �|@      R@     �@     �l@     ȉ@     �u@      <@       @      `@      s@      $@      >@     �i@      =@     ��@     �T@     X�@     `d@      &@              4@     �S@       @      @     �I@             Pq@      9@     �a@      =@      �?              "@      =@               @      3@             �`@      @     �F@       @      �?              @      ,@                      &@              =@      @      (@      @                      @      .@               @       @             �Z@      �?     �@@       @      �?              &@      I@       @      @      @@             �a@      5@     @X@      5@                      @      9@       @      @      6@             @Q@      ,@     �D@      $@                      @      9@               @      $@             @R@      @      L@      &@               @     @[@      l@       @      7@      c@      =@     �y@      M@     �w@     �`@      $@      @     �N@     `a@      @      "@      R@      3@      l@      =@     �n@     @Q@      @      @      =@      I@      @      @     �B@      &@     �I@      ,@     �H@      A@      @              @@     @V@       @      @     �A@       @     �e@      .@     �h@     �A@              @      H@     �U@      @      ,@     @T@      $@     `g@      =@     �`@     @P@      @              0@      :@              @      1@      �?     @W@      @     �I@       @              @      @@      N@      @      &@      P@      "@     �W@      :@      U@     �L@      @      "@      g@     @m@      ,@     �B@     �o@     �E@     s@     `b@     �r@     @g@      1@       @     �C@     @R@      �?       @     �J@      @     @[@      3@     �[@      B@      @       @      <@      N@      �?      @     �D@      @      X@      @     @X@      2@      �?       @      0@      ?@      �?      @      5@       @      L@      @      D@      (@                      (@      =@                      4@       @      D@      �?     �L@      @      �?              &@      *@              @      (@      �?      *@      (@      ,@      2@       @              &@      &@              @      @              @      @      @      *@                               @                      @      �?      "@      @      "@      @       @      @      b@      d@      *@      =@      i@      C@     �h@      `@     �g@     �b@      ,@      @     @Z@     �\@      $@      7@      a@      A@     �S@     �[@     �W@     �]@      ,@      @     @Y@     �\@      $@      7@      `@     �@@     �S@     �X@     @V@      ]@       @              @      �?                       @      �?              &@      @       @      @      �?      D@      G@      @      @      P@      @     @]@      2@     @X@      @@              �?     �@@     �F@       @      @      N@       @     @]@      2@     @X@      @@                      @      �?      �?              @       @                                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ J6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?	��dI@�	           ��@       	                   �;@��'��'	@�           ��@                          �1@}���N�@;           @�@                            �?���{�1@c            �b@������������������������       ����[E@5            �S@������������������������       �:k�h�z@.             R@                           �?{��;�@�           �@������������������������       �`�o$S�@           �|@������������������������       �2qF�	@�           ��@
                          �=@�x���	@�            `q@                           �?��ژ�@L            �^@������������������������       �ࠃ�c@             B@������������������������       ���
�\Z@6            �U@                           �?�x7\�@\            �c@������������������������       �]�f��Y@            �D@������������������������       �{��FQ�@D            �\@                           �?^6���$@�           F�@                           �?���.��@�           ��@                          �6@�Mfo� @	           @y@������������������������       �,����?�            �s@������������������������       ���.�@>            �V@                          �7@�f$MY�@�            �s@������������������������       �Գ��@�            �o@������������������������       �摽 ��@(             P@                           �?�#�.@�           @�@                          �8@\�����@9            �Y@������������������������       ���A�q�@0            �T@������������������������       ���}��9@	             4@                          �4@d��nO�@�           ��@������������������������       �����-�@�           ��@������������������������       ���i!�@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@      s@     0�@      @@      K@     @}@     @R@     `�@     �l@     @�@     �w@     �@@      &@     �d@      m@      7@      >@     �l@      C@     �l@     �c@      n@      h@      7@       @     �`@     `i@      0@      5@     @h@      4@     `k@     �_@      k@     �]@      4@      �?      (@      5@      �?              4@              L@      @      ;@      "@              �?      @      ,@                      $@              3@      @      4@      @                      @      @      �?              $@             �B@      �?      @       @              @     @^@     �f@      .@      5@     �e@      4@     `d@     �^@     �g@     �[@      4@              9@      U@              @     �R@      @      X@      F@     �R@      F@      @      @      X@     �X@      .@      ,@      Y@      0@     �P@     �S@      ]@     �P@      0@      @      ?@      >@      @      "@     �A@      2@      (@     �@@      8@     @R@      @      @      $@      *@      @      @      @      *@       @      (@      0@     �C@      �?      �?      @      @                       @       @                      @      *@               @      @      @      @      @      @      &@       @      (@      &@      :@      �?              5@      1@      @      @      <@      @      $@      5@       @      A@       @              @      @       @               @      �?      @      @      @      $@                      .@      *@       @      @      :@      @      @      0@      @      8@       @      �?     �a@     �q@      "@      8@     �m@     �A@     (�@     �Q@     ��@      g@      $@              <@     @Q@      �?      �?     �H@      @     �t@      $@     �g@      A@      @              ,@      C@              �?      @@      @      j@      @      U@      2@                      @      @@              �?      :@       @     @f@       @     �L@      "@                      @      @                      @       @      >@      @      ;@      "@                      ,@      ?@      �?              1@      @     @^@      @     @Z@      0@      @              (@      ;@      �?               @             @[@      @     �T@       @      @               @      @                      "@      @      (@      �?      7@       @       @      �?     �\@      k@       @      7@     �g@      <@     �{@      N@     �w@     �b@      @      �?       @      .@              $@      .@      @      *@       @      3@      @              �?      @      .@              @      ,@      @      &@      @      2@      @                      @                      @      �?               @      @      �?       @                     �Z@      i@       @      *@     �e@      6@     �z@      J@     pv@     �a@      @             �B@     �Z@      @      @      K@      �?     r@      9@     �e@      M@                     @Q@     �W@      @      @     @^@      5@     �a@      ;@      g@     @U@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @v�[^?@�	           ��@       	                   �4@�h��@�           �@                          �0@�9�m�@d           ��@                            �?��w�R�@e             c@������������������������       ���_-!��?!             K@������������������������       ������ @D            �X@                           �?S_����@�           $�@������������������������       �q([Wyr@           �y@������������������������       �)՜���@�           ��@
                           @�4�`l@�           ��@                           �?&і¢	@�           ��@������������������������       ��.B�	@g           �@������������������������       �Ȭ�}$@�            �j@                          �7@���g�@�           `�@������������������������       ��&Sx2@�            ps@������������������������       �
��Aٷ@�            Pu@                           @+,����@�           �@                           �?=>~켟@            �@                          �8@#W`@�            �m@������������������������       �><�v��@u            `f@������������������������       ��8t*{A@&            �L@                          �?@����:	@{           ��@������������������������       ����i�@i           ؁@������������������������       �%�xi�@             =@                          �=@��� �)@�            0p@                           �?�	dy�@�            �m@������������������������       �;/��)�?:             X@������������������������       ��=a�s�@f            �a@������������������������       �L�� @	             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �q@     Ѐ@      5@      N@     �z@     @X@     D�@     �l@     �@     �w@      ;@      @     @i@     Px@      .@     �B@     `q@     @Q@     ��@     �d@     8�@     pp@      8@      �?      P@     �e@      �?      $@     @]@      ,@     `@     �Q@     @r@     �^@       @                     �C@                      $@              K@       @      ;@      4@                              &@                       @              9@       @      �?      *@                              <@                       @              =@              :@      @              �?      P@     �`@      �?      $@     �Z@      ,@      |@     @Q@     �p@     �Y@       @              4@     �E@              @      1@      �?     `f@      2@     �Y@      9@      �?      �?      F@      W@      �?      @     �V@      *@     �p@     �I@     `d@     �S@      @      @     @a@     �j@      ,@      ;@      d@     �K@     �q@     �W@     0r@     �a@      0@      @     @X@     @Z@      $@      6@     �X@     �B@     �Y@      Q@      `@     �Y@      *@      @     �Q@      S@      $@      2@      T@      9@      Q@     �G@     @T@     �U@      $@              ;@      =@              @      2@      (@     �A@      5@      H@      .@      @             �D@     �[@      @      @     �O@      2@     �f@      ;@     @d@      C@      @              2@      O@       @      �?      7@       @      \@      @     �P@      $@       @              7@      H@       @      @      D@      $@     @Q@      5@     �W@      <@      �?      (@     �S@     �b@      @      7@     �b@      <@     �o@      O@     �j@     @\@      @      (@     �Q@      `@      @      3@     �`@      ;@     �c@      M@      `@      W@      @              6@      A@      �?      @      6@              Q@      (@     �G@      7@                      (@      8@      �?      �?      ,@              M@      @     �E@      3@                      $@      $@              @       @              $@      @      @      @              (@      H@     �W@      @      (@     @\@      ;@      V@      G@     �T@     @Q@      @      @     �D@     @W@      @      &@     @Z@      ;@      V@     �F@      T@     �P@      @      @      @       @              �?       @                      �?       @       @                      "@      4@              @      0@      �?     �X@      @     @U@      5@                      "@      3@              @      ,@      �?      X@      @     �S@      *@                      @      @              �?      @              J@      @      =@                              @      0@              @      &@      �?      F@      �?      I@      *@                              �?                       @              @              @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ"��[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Uɥi��@�	           ��@       	                    �?D��4kI@           H�@                          �3@I�$ه@B           �~@                           �?Af�r�P@s            �d@������������������������       ��(o��@0             Q@������������������������       �Hz�^NB@C            �X@                            �?�\յ��@�            `t@������������������������       ��7Ρl@q             e@������������������������       �A ���@^            �c@
                           �?�i��z�@�           (�@                            �?�
�R � @�            0x@������������������������       ���/^l�?:            �W@������������������������       ���5^�Q@�            Pr@                           @IH�j@�             v@������������������������       ���0h�@�            @h@������������������������       �5�kE�@X             d@                            @�;���@�           �@                          �;@����:N@�           p�@                           @���{�@           ,�@������������������������       �)��*}@|           (�@������������������������       ��H�Ȃ�@�           �@                          �?@D��y��@�             j@������������������������       ��*�Y�N@j            �d@������������������������       ��P}v@            �E@                           �?����@�           ؈@                           �?a���~B@8            �V@������������������������       ��A;@&            �N@������������������������       �)���@             >@                           �?U����@�            �@������������������������       �J\6 �	@           �z@������������������������       �	3��{@�            @q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@     �@      6@     �K@     �z@     �V@     �@     �i@     0�@     `w@      5@      �?     @W@     �b@       @      "@     @]@      @     `|@     �A@     �q@     @S@      @      �?     �L@     �P@      �?       @      Q@             �Z@      ;@     �[@     �F@       @              "@      3@               @      4@              I@      (@      A@      5@                               @                      "@              7@      @      2@      @                      "@      &@               @      &@              ;@      "@      0@      ,@              �?      H@      H@      �?      @      H@             �L@      .@      S@      8@       @      �?      ?@      1@      �?       @      1@              ;@      @     �G@      1@       @              1@      ?@              @      ?@              >@      "@      =@      @                      B@     �T@      �?      �?     �H@      @     �u@       @     �e@      @@      @              6@      D@              �?      7@      @     �i@      @     @R@      0@                              @              �?      @      �?     �N@              0@      @                      6@      B@                      1@       @      b@      @     �L@      &@                      ,@      E@      �?              :@      @     �a@      @     �Y@      0@      @              $@      7@                      "@      @      U@             �J@      "@       @              @      3@      �?              1@              M@      @     �H@      @      �?      .@     �i@     �v@      4@      G@     �s@     �T@     ��@      e@     H�@     �r@      0@      @     `a@      p@      &@      ;@      l@     �H@      ~@     �]@     pw@     �g@      "@      �?     �_@      m@       @      :@     `f@      ?@     �|@     �Y@     Pu@     �c@       @             �Q@      b@      @      .@     @^@      9@     �q@      D@     �k@     �Z@      @      �?     �K@      V@      @      &@      M@      @     �f@      O@     �]@     �J@      @      @      *@      7@      @      �?     �F@      2@      3@      1@      A@      ?@      �?      @      @      ,@      @      �?     �D@      ,@      ,@      1@      @@      4@      �?               @      "@                      @      @      @               @      &@              $@     �P@     �[@      "@      3@      V@      A@     �b@      I@     @b@     �Z@      @       @      ,@      0@              @      ,@      @      @      0@      (@      @               @       @       @                      *@      @      �?      *@      &@      �?                      @       @              @      �?       @       @      @      �?      @               @     �J@     �W@      "@      0@     �R@      <@      b@      A@     �`@     �Y@      @       @     �E@      K@       @      $@     �J@      :@      L@      8@     �P@     @R@      @              $@      D@      �?      @      5@       @     @V@      $@     �P@      =@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ%O`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�t�t]@�	           ��@       	                    �?G��o�@z           ~�@                           �?~=���4	@           ��@                           �?�Su@�           �@������������������������       ���W
_D@u            �h@������������������������       ��gkR@           �y@                          �8@�:L##�	@�           p�@������������������������       ���_�I	@�           H�@������������������������       �p�r�+�	@�            0u@
                            �?5�-���@g            �@                          �1@���Ի@�            pu@������������������������       �n��[�>@             �N@������������������������       ��Ӻ.�7@�            �q@                            @2�oY�7@�             m@������������������������       ��&L��W@7             U@������������������������       �ѳ]��@_            �b@                          �4@�0�E@5           (�@                           �?�-�ZZ@O           ��@                          �1@~|���?�            �t@������������������������       �����"��?Z            @`@������������������������       ���؆��?�            �i@                          �1@��%ʞ�@m           8�@������������������������       �����#z @�             i@������������������������       �u�`�v=@�            �w@                           @�ԕ���@�           ��@                          �5@�R�D6�@6           �~@������������������������       ���Y�5�@E            @\@������������������������       �MN���@�            �w@                           �?�[�m��@�            `p@������������������������       �`d�7@U             a@������������������������       ���C�"(@[            @_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     h�@      >@     �C@     �|@      V@     x�@      l@     @�@     �v@      ;@      8@      m@     �t@      6@      ;@     �s@     �Q@     �w@     �g@     px@     `m@      4@      8@     �f@     �m@      4@      8@     �n@      L@     @n@     �b@     `q@     �g@      3@      @     �H@      X@       @      $@     @W@      "@      a@      B@     �Z@     @P@      @       @      8@      ;@                      9@              M@       @      I@      "@      �?      �?      9@     @Q@       @      $@      Q@      "@     �S@      A@     �L@      L@      @      5@     �`@     �a@      2@      ,@      c@     �G@     @Z@      \@     `e@      _@      .@      0@     �U@      X@      &@       @     �]@      9@     �T@      M@     �`@     �P@      $@      @     �F@      F@      @      @      A@      6@      7@      K@      B@      M@      @             �I@     @X@       @      @     �Q@      ,@      a@     �E@     @\@      G@      �?              B@      N@       @      @      B@      "@     �R@      2@     @T@      7@      �?              @      $@                      �?              <@      �?      &@      @                      =@      I@       @      @     �A@      "@      G@      1@     �Q@      4@      �?              .@     �B@                      A@      @      O@      9@      @@      7@                      @      @                      5@       @      2@      &@      1@      @                      (@      >@                      *@      @      F@      ,@      .@      2@              �?     @U@      l@       @      (@     �a@      2@     ��@     �@@     z@     @`@      @              >@     �Z@      @      @     �G@      @     `y@      1@     �l@     �M@      @              @      ;@               @      $@              i@       @     @R@      $@      @                      &@              �?       @             �T@              9@              @              @      0@              �?       @             �]@       @      H@      $@                      7@      T@      @      @     �B@      @     �i@      .@     �c@     �H@                      @      =@               @      @             @U@       @     �O@      $@                      4@     �I@      @      @      >@      @     @^@      *@     �W@     �C@              �?     �K@     @]@      @      @     �W@      (@     �g@      0@     `g@     �Q@      @      �?     �E@     �P@              �?     �M@      @     @b@      @     @^@      E@      @              @      6@                      2@      �?      <@      �?      A@      @      @      �?      D@     �F@              �?     �D@      @     �]@      @     �U@     �C@      �?              (@      I@      @      @      B@      @     �F@      &@     �P@      =@                      @      =@              @      6@       @      5@       @     �C@      *@                      @      5@      @              ,@      @      8@      "@      ;@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@����Dg@�	           ��@       	                    @+T��ۯ@�           D�@                           @%���ޮ@�           Є@                           �?�č��@           �{@������������������������       �l6�~Pk@c            �a@������������������������       �C7V�R�@�            �r@                           @��j>�D@�             l@������������������������       �Vz�+s@~            �g@������������������������       �,�|#��@            �A@
                           �?�/��@�           ��@                          �0@��TM�Y�?�            s@������������������������       ��ߘ�G`�?+            @Q@������������������������       ��s\Y�?�            �m@                           @����-@           `|@������������������������       ���R=�@?            �[@������������������������       �����"@�            �u@                           �?U��	�@!           p�@                           @h�N���@�           �@                          �<@��3m�@           �z@������������������������       �ɯ{�^@�            Pv@������������������������       �R\e�t=@,            @Q@                          �>@q��]V�@�            0q@������������������������       �fLu	@�            �p@������������������������       �lofON@             &@                           @R~��{,	@a           �@                          �9@>7���	@�           ܐ@������������������������       ��[���	@�           ��@������������������������       ��U��E
@�             v@                          �7@��[�5@�            �@������������������������       �i<�)�.@           Py@������������������������       ��P"%�,@�            �r@�t�b�N      h�h5h8K ��h:��R�(KKKK��h��B�        2@     r@     8�@      @@      J@     �{@     �X@     0�@      l@      �@     `u@      A@       @     �S@     �g@      @      @     ``@       @     @      P@     t@     �]@      @       @     �G@     �W@      @      @     �S@      @     @d@      I@     `a@     @S@      @      �?     �B@     �N@       @      @      I@      �?      [@      7@     �[@      F@              �?      $@      5@      �?              8@             �D@      &@      :@      @                      ;@      D@      �?      @      :@      �?     �P@      (@     @U@     �B@              �?      $@      A@      �?              =@      @      K@      ;@      <@     �@@      @              $@      =@      �?              6@      �?      I@      7@      8@      <@       @      �?              @                      @      @      @      @      @      @      �?              @@      X@       @       @      J@       @     �t@      ,@     �f@     �D@      �?              &@      >@              �?      "@             @e@       @      P@      &@      �?                      ,@                      @             �A@              &@      @                      &@      0@              �?      @             �`@       @     �J@      @      �?              5@     �P@       @      �?     �E@       @     �d@      @     �]@      >@                      (@      <@                      @       @      C@       @      (@      &@                      "@      C@       @      �?      C@             �_@      @     �Z@      3@              0@     @j@     �x@      ;@     �G@     ps@     �V@     P@      d@     �}@      l@      >@      �?      O@     �_@      �?      @     �N@      "@     `j@      <@      a@     �J@      @      �?     �J@      S@              @     �F@       @     @X@      6@      S@      E@      @      �?      G@      N@              @     �@@       @     @W@      0@      R@      9@      @              @      0@               @      (@              @      @      @      1@      �?              "@      I@      �?              0@      @     �\@      @     �N@      &@                      "@     �H@      �?              *@      @     @\@      @      N@       @                              �?                      @              �?       @      �?      @              .@     �b@     �p@      :@      D@     @o@     @T@      r@     �`@     `u@     `e@      9@      ,@     �Z@     �f@      5@     �@@     @f@      O@     �W@      Y@     �b@     �^@      2@      "@     �P@     @`@      *@      <@      a@      =@     �P@     �K@     �Z@     @S@      $@      @      D@     �I@       @      @     �D@     �@@      <@     �F@     �E@     �F@       @      �?      E@     @U@      @      @      R@      3@     �h@     �@@      h@     �H@      @              2@      N@      @      @      ;@      0@      `@      @     �\@      3@      @      �?      8@      9@              �?     �F@      @      Q@      ;@     �S@      >@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJWG�]hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �8@�e�^@�	           ��@       	                    @[��Q@R           �@                           �?�����@�           ��@                           �?�%e�[@D           �@������������������������       �<�W�5@�            Pv@������������������������       �wv���@b            �b@                          �3@a���y�@�           ��@������������������������       �*Y5L�@           �z@������������������������       �'�p��@�           ؃@
                          �4@����@n           ��@                           @�=e�o�@H           ��@������������������������       � ��0��@�            �j@������������������������       �=���<@�           ��@                           @^$ʹ��@&           �}@������������������������       ��C�0�@F            @[@������������������������       �=��Ѷ@�            �v@                           �?��Tw��	@S           ��@                           �?��-kP
@A           p�@                           �?�v�Q��@M            �[@������������������������       ��bn�@             �D@������������������������       ���y	A$@-            @Q@                          �;@d5�U
@�             z@������������������������       ��l��/�	@s            �f@������������������������       �UI?�k�	@�             m@                           @�gAOc�@           �z@                           �?q~۪��@           Py@������������������������       �~<�\��@I            �Z@������������������������       �8�Ə��@�            �r@������������������������       �Q�	�n@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        5@     �s@     ��@     �@@      L@     `|@      S@     ��@     `m@     H�@     �u@     �E@      $@     �k@     �x@      8@      @@     �u@     �D@      �@     �_@     x�@     `j@      7@      $@     �b@     �k@      1@      6@     �n@      >@      t@      [@     �q@     `b@      *@             �I@     @P@      @      @      K@      �?     �c@      8@     �\@      >@      @             �A@      K@      @      �?     �D@      �?     �V@      6@     �S@      ;@      @              0@      &@               @      *@             @P@       @      B@      @              $@     @X@     �c@      ,@      3@      h@      =@     �d@      U@     @e@     @]@      $@      @      :@     �N@      �?       @      L@      *@     �W@      B@     �R@      K@      @      @     �Q@      X@      *@      1@      a@      0@     �Q@      H@     �W@     �O@      @             �R@     �e@      @      $@     �Y@      &@      �@      3@      u@      P@      $@              E@     �X@      @      "@      L@       @     �z@      $@     �k@      D@      @              3@     �C@                      &@       @     �U@      @     �F@      "@                      7@     �M@      @      "@     �F@             `u@      @     @f@      ?@      @              @@      S@       @      �?      G@      "@      c@      "@     �\@      8@      @              "@      5@                      @      @      D@              4@      @      @              7@     �K@       @      �?     �C@      @      \@      "@     �W@      5@      @      &@     @X@     �`@      "@      8@     �Z@     �A@     �^@      [@     @c@     @a@      4@      &@     �N@     �V@      @      (@      J@      6@      D@      N@      N@     �V@      3@              (@      9@              @      $@      �?      .@      @      2@      3@                      @      @                      @              @      �?      @      $@                      @      2@              @      @      �?       @      @      (@      "@              &@     �H@     �P@      @      "@      E@      5@      9@     �J@      E@      R@      3@      �?      3@      <@      @      @      3@      $@      0@      A@      :@      .@      "@      $@      >@      C@      @      @      7@      &@      "@      3@      0@     �L@      $@              B@     �D@       @      (@      K@      *@     �T@      H@     �W@     �G@      �?              ;@     �D@       @      (@     �H@       @     @T@     �F@      W@     �G@      �?              @      @                      "@      @      @@      $@      ?@      &@      �?              8@      B@       @      (@      D@      @     �H@     �A@     �N@      B@                      "@                              @      @      �?      @       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Z�DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @����b@�	           ��@       	                   �4@�	<� @�           ��@                           �?�l��@C           |�@                           @fҮRZ�@,           �}@������������������������       �{})��@z             j@������������������������       ���x-�L�?�            �p@                           @�Q0�2c@           �@������������������������       �}�|�s@�            �t@������������������������       �VB��@3           �@
                           @�Mw��e@�           ̖@                           �?��>5��@5           0�@������������������������       ��� ��_	@W           h�@������������������������       �n.�|R�@�           ��@                           @���-	@h            �d@������������������������       �
��$\�	@C            �[@������������������������       �V�x@��@%            �L@                           �?�7M�� @�           ܑ@                          �>@�)�=�@�             t@                           �?z����@�            @s@������������������������       �,<��"@q            @g@������������������������       �ُ�I�D�?[            �^@������������������������       ��bN�� @             ,@                           �?$\��C�@�           ��@                           �?����@*             S@������������������������       �4l ��?             4@������������������������       �~=&υ�@             L@                           �?�֭@j@�           H�@������������������������       �X�y�@�            �q@������������������������       ���<�8�@           �|@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     �q@      �@      ?@     �L@     �~@     �U@     ��@      j@     �@      v@      >@      $@     �g@     �z@      .@     �B@     @t@     �P@     ؅@     `a@     �@     �m@      3@             �Q@     @g@      @      $@      _@      @      |@      M@     �r@     �Y@      @              :@      J@              �?      F@      �?     �i@      (@      [@      :@       @              (@      8@                      =@      �?      K@      "@      M@      3@       @              ,@      <@              �?      .@             �b@      @      I@      @                      F@     �`@      @      "@      T@      @     �n@      G@     �g@     @S@      �?              <@      N@       @      @     �G@      @      N@      B@     �H@     �C@      �?              0@     �R@       @      @     �@@             @g@      $@     �a@      C@              $@     @^@     �m@      &@      ;@      i@      O@      o@     @T@     `s@     �`@      0@      @     �X@     �k@      @      ;@     �e@      J@     @m@      H@      r@     �^@      *@      @      N@     �W@      @      1@     �V@      ;@      G@      ?@     �S@     �N@      @      �?     �C@     �_@      �?      $@     �T@      9@     �g@      1@     `j@     �N@      @      @      6@      1@      @              <@      $@      .@     �@@      4@      (@      @      @      .@      *@      @              (@      "@      @      9@      $@      "@      @              @      @                      0@      �?       @       @      $@      @              @     �V@      g@      0@      4@     �d@      5@     �n@     @Q@      h@     @]@      &@              :@      H@      �?      @      B@      �?     �[@      .@      P@      0@                      :@      H@      �?      @      >@      �?     �[@      *@     �N@      .@                      4@     �F@      �?      @      6@      �?      G@      (@      9@      &@                      @      @                       @              P@      �?      B@      @                                               @      @                       @      @      �?              @     @P@      a@      .@      .@     ``@      4@      a@      K@      `@     @Y@      &@      @      @      5@              @      &@      @              ,@      @      @              �?              *@                              @              @                              @      @       @              @      &@       @              &@      @      @              @      M@     �\@      .@      &@      ^@      .@      a@      D@     �_@     �W@      &@       @      2@      F@      &@      @     �G@       @      E@      *@      K@      C@       @      �?      D@     �Q@      @      @     @R@      @     �W@      ;@      R@      L@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��4`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�J��!@�	           ��@       	                   �5@ZH���@           T�@                           @:�z@�#@�            �@                          �1@�"��
�@�            �v@������������������������       �h�$,�@C             \@������������������������       �wtq�4D@�            �o@                           @�v�!i�?�            Py@������������������������       ��&��Y��?�            �q@������������������������       ��?Ѥ@M             _@
                          �=@����`!@2           }@                          �<@RB2��\@
           py@������������������������       � ���3@�            Pw@������������������������       ������@             A@                            �?�t��T�@(             M@������������������������       �����@	             1@������������������������       ��"�a׹@            �D@                           @PŌ��!@�           �@                           �?8��ˊ	@�           |�@                           @2�}*��	@�            �@������������������������       ����w-�	@�           ��@������������������������       �-��O�	@�            �v@                           �?ȯ�@           �y@������������������������       ���F��-@             <@������������������������       ���h�ȧ@�            0x@                           @t����@�           T�@                           @��c�3@�           $�@������������������������       ���^"�d@�           (�@������������������������       ��h��Y�@�            @r@                          �4@��XHI@U            �a@������������������������       ��(��� @            �K@������������������������       �7�R`X`@6            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     @r@     P�@      4@     �G@      |@     �T@     ��@     �i@     �@     �w@     �C@             @R@     �b@       @      &@     �X@      @     �}@     �C@     �q@      V@      @             �@@      V@              @      D@      @     �v@      1@      e@      H@      @              4@      B@              @      >@      @     @_@      ,@     @V@     �D@      �?              @      *@                      .@              E@      @      ;@      @                      ,@      7@              @      .@      @     �T@      $@      O@      B@      �?              *@      J@                      $@             �m@      @      T@      @       @              $@      @@                      @             `f@             �J@      @                      @      4@                      @             �M@      @      ;@      @       @              D@     �O@       @      @     �M@       @      ]@      6@     @\@      D@      @             �A@     �L@       @       @      H@      �?     @[@      3@     @Y@     �@@                      =@      I@       @       @     �G@      �?      Y@      2@     �X@      :@                      @      @                      �?              "@      �?      @      @                      @      @              @      &@      �?      @      @      (@      @      @               @      �?                      @      �?                      �?      @      @              @      @              @      @              @      @      &@      @              4@     `k@     0w@      2@      B@     �u@      S@     (�@     �d@     �@      r@     �@@      2@     `d@      j@      1@      9@     `m@      P@     `h@      a@     �k@     @h@      <@      2@     �_@      b@      .@      2@     �f@     �H@     �^@     @W@     �a@     �b@      ;@      *@      U@      U@      &@      @     @`@      E@      S@      L@      Z@     �Y@      *@      @      E@     �N@      @      &@      J@      @     �G@     �B@     �C@     �G@      ,@             �B@     �O@       @      @     �J@      .@      R@     �E@     @S@     �F@      �?              @       @              @      @                       @       @      @                      @@     �N@       @       @      G@      .@      R@     �D@     �R@      D@      �?       @      L@     `d@      �?      &@      ]@      (@      x@      >@     pr@      X@      @       @     �E@     �b@      �?      "@      Z@      $@     �t@      6@     0q@      U@               @      ?@     �[@              @     �R@      @      p@      (@     �h@      G@                      (@     �B@      �?      @      =@      @     @S@      $@     @S@      C@                      *@      .@               @      (@       @     �I@       @      4@      (@      @              @      @               @                      =@       @       @      @                      "@      (@                      (@       @      6@      @      (@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ;�KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?c���sk@�	           ��@       	                    @�"$z=�@           X�@                           �?<;��<�@�           p�@                           �?��"��@             i@������������������������       �/q�+�r@>            @X@������������������������       ��{i��B@A            �Y@                            �?��1�8S@'           `|@������������������������       ����ڦ�@Q            @^@������������������������       �|�Kӟ@�            �t@
                           �?��&}V� @k           @�@                          �;@h���'@�            @v@������������������������       �����@�            �t@������������������������       � ��$���?             7@                           @���st/ @�            �l@������������������������       ��ƴ=���?N             _@������������������������       ��wf�% @D             Z@                          �4@o��J@�           �@                          �1@�0p5x@�           ,�@                           �?�`����@�            �v@������������������������       �q�t�(@:            �V@������������������������       ��F����@�            Pq@                           �?��Å_@�           ��@������������������������       �Ɯ&�@#            �N@������������������������       ����^\@�           ��@                          �:@�^�	@�           ��@                          �7@�*J{@�           ��@������������������������       ��Nz�@�           p�@������������������������       ��Z��n�@            {@                          �<@�]W�	@           �z@������������������������       ��}��	@{            �f@������������������������       ����K�@�            `n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     `u@     ��@      ;@      K@     P|@     @U@      �@     `k@     �@      v@     �B@      @      T@     �d@       @      $@     @Z@      $@     �{@      E@     �q@     �T@      $@      @      O@     @U@      �?      "@     @R@      @     �c@     �B@      c@      N@      "@      @      $@      @@                      7@              M@      @     �J@      ,@      @      @      @      0@                      "@              =@      @      :@      @                      @      0@                      ,@              =@      �?      ;@      "@      @              J@     �J@      �?      "@      I@      @      Y@     �@@      Y@      G@      @               @      3@               @      "@      �?      :@      @      D@       @       @              F@      A@      �?      @     �D@      @     �R@      ;@      N@      C@      @              2@     �S@      �?      �?      @@      @     r@      @     @`@      6@      �?              *@     �I@              �?      9@      @     @f@      @     �P@      ,@                      *@      G@              �?      9@      �?     �d@      @     �P@      ,@                              @                              @      ,@              �?                              @      <@      �?              @       @     �[@       @     �O@       @      �?              @      "@                      �?       @     �Q@      �?     �A@       @                       @      3@      �?              @              D@      �?      <@      @      �?      ,@     `p@      w@      9@      F@     �u@     �R@     �@      f@     @�@     �p@      ;@       @     �S@     �b@       @      .@     �a@      .@     @u@      P@      o@     �U@      $@      �?      3@     �G@      �?      @     �A@      �?     �a@      &@      V@      .@              �?      $@      "@      �?      @      0@      �?      4@      �?      8@      @                      "@      C@               @      3@             �^@      $@      P@      (@              �?      N@      Z@      @      "@      [@      ,@     �h@     �J@      d@      R@      $@               @      @              �?      *@      �?      @       @      5@      @              �?      M@     @X@      @       @     �W@      *@      h@     �F@     �a@     @Q@      $@      (@     �f@      k@      1@      =@     �i@      N@     �i@     @\@     �p@     �f@      1@      @      ^@     @f@      @      6@      b@     �B@      d@     �S@     �k@     @Y@      *@      @     @W@      ]@      @      0@      U@      2@     @W@     �A@     �`@     �J@      @              ;@      O@      @      @      N@      3@      Q@     �E@     �U@      H@       @      "@     �O@     �C@      $@      @     �N@      7@      F@     �A@     �H@     �T@      @      @      8@      (@      @      @      5@      @      =@      1@      :@      >@      @       @     �C@      ;@      @      @      D@      2@      .@      2@      7@      J@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�9HhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Z���R@�	           ��@       	                   �8@J�0��@t           �@                           �?�A�(�1@�           h�@                           �?2��Ζ@�           8�@������������������������       �;��%*m@�            �u@������������������������       ��TUC	@�           ��@                           �?%xW�Ñ@.           �|@������������������������       ����j@Z            �b@������������������������       �MU���@�            �s@
                           �?��	@�           8�@                          �;@(1���	@7            ~@������������������������       ���m�	@�            �m@������������������������       ���Ne��@�            �n@                           @���;v@R            �`@������������������������       ��,z�#B@;            �W@������������������������       ����"@            �C@                           �?��冽�@J            �@                          �3@&�ġ� @o           ��@                           @�XM��
�?�            �s@������������������������       �39��ه�?+            �Q@������������������������       �H�Vw*��?�             o@                            @��G!­@�            Pq@������������������������       �ܕ��@�            �l@������������������������       �,�gp�)�?            �H@                           @Q/�@�           Б@                           @%v>���@�           `�@������������������������       �wc �U@�           h�@������������������������       ��j��@�            �t@                          �:@�?�:@             <@������������������������       �g�n�	@             2@������������������������       ���&��?             $@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     pq@     X�@      >@      K@     �|@     �T@     �@     `n@     �@     �v@     �A@      &@     �h@     �t@      7@      C@     0t@     @P@     �s@     �i@     Px@     �n@      >@      @     �a@      m@      *@      ;@      n@     �E@     pp@     �\@     �s@     `b@      ,@      @      [@     @f@      $@      3@      f@     �@@     �b@      W@     �i@     @]@      (@              ;@      Q@               @     �D@      @      P@      ,@      V@      >@      @      @     @T@     �[@      $@      &@      a@      >@      U@     �S@      ]@     �U@      "@             �A@     �K@      @       @      P@      $@     �\@      7@     �\@      >@       @              ,@      @              �?      ,@      �?      N@       @     �D@       @                      5@      H@      @      @      I@      "@     �K@      5@     �R@      6@       @      @      L@     @X@      $@      &@     �T@      6@      J@      W@     �Q@      Y@      0@      @     �D@     �R@      $@       @     �O@      5@      @@     @R@     �J@     �T@      0@      �?      2@      B@      @      @     �A@      $@      7@     �D@      ?@      4@      $@      @      7@     �C@      @      @      <@      &@      "@      @@      6@     �O@      @              .@      6@              @      3@      �?      4@      3@      1@      1@                       @      0@              @      3@      �?      (@      .@      @      *@                      @      @                                       @      @      $@      @                      T@      l@      @      0@     �a@      1@     0�@      B@     �y@     �]@      @              4@      Q@      �?      @      =@       @     0s@       @     �`@      8@                      "@     �A@              �?      @             �f@       @     @S@      @                              .@                                     �B@              0@       @                      "@      4@              �?      @              b@       @     �N@      @                      &@     �@@      �?       @      7@       @     @_@      @     �L@      1@                      &@     �@@      �?              4@       @     �W@      @     �G@      ,@                                               @      @              >@      �?      $@      @                      N@     �c@      @      *@     �[@      .@     0w@      <@     �q@     �W@      @             �J@     `c@      @      (@      Z@      &@      w@      ;@     `q@     @W@      @              A@     �Z@              @      P@      @     �q@      2@     �i@     �K@      �?              3@      H@      @      @      D@      @      U@      "@     �Q@      C@      @              @       @       @      �?      @      @      �?      �?       @      �?                      �?       @       @      �?      @      @      �?      �?       @      �?                      @                              @                                                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>ޓbhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�ɂ�s&@�	           ��@       	                   �1@I/�nup@Y           ��@                          �0@��s�M@�           x�@                           @� �	��@|            �i@������������������������       ��Q>܋]@f             d@������������������������       �����h��?             F@                           �?���	}@            z@������������������������       �@fU�Z@N             `@������������������������       ��j\�� @�             r@
                           �?�i�G@�           8�@                          �3@�DP:�?@:           P�@������������������������       �1A9S^@�            �r@������������������������       ��-��v�@�            �k@                            �?��m��@�           �@������������������������       ��C�P�@�            0p@������������������������       ���&}�W@�           �@                           �?I���@V           0�@                          �;@\8��c	@"           h�@                           �?Z�
��@{           �@������������������������       �I��E��@g            �d@������������������������       �)/13�z	@           �{@                          �=@O�ǋAS	@�             q@������������������������       ��	���@O             _@������������������������       �_�lTf�@X            �b@                           @4�x�e�@4           ��@                           �?��C�@�            �p@������������������������       �Apw��{@-            �S@������������������������       �"��y@y            �g@                          �7@�+V��@�           ��@������������������������       ��ysuW@�             i@������������������������       �k�v
@           �x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     q@     ��@      :@      G@     @~@      Q@     H�@      j@     ��@     w@     �C@      "@     �Y@     `s@      *@      3@      n@      5@     ��@      V@     �@     �d@      "@      @      :@     �R@      �?      @     �H@      �?     �o@      3@     �b@      F@                      @      B@               @      :@              V@      �?      C@       @                       @      7@               @      :@             �P@      �?      B@      @                      @      *@                                      5@               @      @              @      4@      C@      �?      @      7@      �?     �d@      2@     �[@      B@              @      (@      0@      �?              *@      �?      ;@      @      >@      6@                       @      6@              @      $@              a@      .@     @T@      ,@              @     @S@     �m@      (@      ,@      h@      4@     `{@     @Q@     @v@     @^@      "@              :@     @P@              @     �D@       @     �h@      *@      a@      A@      �?              ,@     �A@              �?      5@             �Z@      (@      V@      8@                      (@      >@              @      4@       @      W@      �?     �H@      $@      �?      @     �I@     `e@      (@      $@     �b@      2@     �m@      L@     `k@     �U@       @              .@     �E@                      H@       @     �P@      5@      F@      2@      �?      @      B@      `@      (@      $@     �Y@      0@     �e@     �A@     �e@     @Q@      @      $@     @e@     �o@      *@      ;@     `n@     �G@     ps@     @^@     ps@     �i@      >@      $@     �Z@     �b@       @      0@      a@      @@     �Q@     �R@     �`@      ]@      8@       @     �U@      Y@      @      @     �Z@      3@      M@      J@     @V@     �N@      4@              <@      >@               @     �@@              3@      @      C@      @       @       @      M@     �Q@      @      @     @R@      3@     �C@     �F@     �I@      L@      2@       @      5@     �H@      @      "@      ?@      *@      *@      6@      F@     �K@      @      @      "@      :@      @      @      ,@      $@      @       @      1@      ;@      @      @      (@      7@              @      1@      @      @      4@      ;@      <@      �?             �O@      Z@      @      &@     �Z@      .@      n@     �G@     @f@      V@      @              9@     �B@              @      B@       @      M@      <@     �E@      8@      @              @       @                      @       @     �@@      @      2@      @      �?              5@     �A@              @      =@      @      9@      7@      9@      2@       @              C@     �P@      @      @     �Q@      @     �f@      3@     �`@      P@      @              (@      @@      @       @      4@       @     �Q@      �?     �E@      .@                      :@     �A@       @      @      I@      @     �[@      2@      W@     �H@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ 3�;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�L���@�	           ��@       	                    �?��̆U�@           ��@                            �?����a@�           H�@                           �?U��!)�@g            �e@������������������������       ��2�3��@'            �P@������������������������       �K��=0�?@            �Z@                          �4@�=R���@-           �@������������������������       �D�SN�� @�            �p@������������������������       ��FQ��@�            �n@
                          �4@�m��g�@q           �@                           �?�f`�E@�            @t@������������������������       �r���@I            �[@������������������������       ���A�r��?{            �j@                            @ɺ���@�            �o@������������������������       ���|R�Y@z            `f@������������������������       ���qA@�@3            �R@                           �?K����@�           ��@                            @�,��z@	@�            @k@                            �?�=���@O            �^@������������������������       ��s��}@?            �W@������������������������       �ޯ5��@             ;@                           �?3�����@4             X@������������������������       ��J��[k@             @@������������������������       �W�ۂ�@#             P@                            @U>�^`�@%           
�@                            �?��o@j           ��@������������������������       �N7�=�@Z           ��@������������������������       �^���@           �z@                          �3@��&��@�           ��@������������������������       ���o+��@�            �k@������������������������       �~��/�	@4            |@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �q@     @@      =@     �P@     `{@      P@     đ@      j@     ��@     �u@      8@              S@      b@      @      &@     @X@      @     (�@      F@     �q@     @S@      @              C@     �Q@      @      @     �K@      @     �r@      <@     �a@      A@      �?                      5@               @      2@      �?     @S@      @      D@      @                              (@              �?      "@      �?      2@      @      1@      �?                              "@              �?      "@             �M@              7@      @                      C@      I@      @      @     �B@      @     �k@      5@      Y@      <@      �?              (@      8@              �?      (@      �?     �a@      "@      K@      @      �?              :@      :@      @       @      9@       @      T@      (@      G@      5@                      C@     @R@              @      E@              k@      0@     �a@     �E@       @              .@      B@              @      1@             �c@      @     �R@      0@                      @      3@              @      $@              ?@      @      ;@      "@                       @      1@                      @             �_@       @     �G@      @                      7@     �B@               @      9@              N@      &@     �P@      ;@       @              0@      5@               @      2@              C@      @      L@      4@       @              @      0@                      @              6@      @      $@      @              :@      j@     @v@      8@     �K@     Pu@      N@     `�@     �d@      �@     �p@      5@      @      ;@      =@               @      A@       @      6@      5@      D@      5@      �?      @      ,@      &@              @      ,@      @      4@      @      >@      (@      �?      @      "@      @              @      (@      �?      0@      @      7@      &@      �?      �?      @      @                       @      @      @              @      �?              @      *@      2@              @      4@      @       @      ,@      $@      "@              @       @      ,@                      @       @              @       @      @                      &@      @              @      1@       @       @      &@       @      @              3@     �f@     pt@      8@     �G@     0s@      J@     ��@     �a@     �}@     �n@      4@      "@     @a@      n@      $@      B@      j@     �B@     |@     @\@     �u@      e@      @      "@     �Z@     @f@      "@     �@@     @b@      >@     pt@     @W@     Pp@     �a@      @              ?@      O@      �?      @     �O@      @     �^@      4@      V@      =@      @      $@     �E@     �U@      ,@      &@     �X@      .@     �b@      >@     �^@     �S@      *@       @       @      >@      �?              A@      @      P@       @      G@      :@               @     �A@     �L@      *@      &@      P@      &@     @U@      6@     @S@      J@      *@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �<@W�l�q@�	           ��@       	                   �3@{Ȼy@�            �@                           �?�O��e@�           ��@                          �2@�,�V�k@g           p�@������������������������       ���c�@           �z@������������������������       ��!��@U             `@                          �1@�ׇy��@)           ��@������������������������       ��z���@�            �t@������������������������       �_\�-wR@S           p�@
                           @Y��[�@J           ��@                           �??�Ay~�@           ��@������������������������       ��@�Æ�@�            �v@������������������������       �,���)	@=           ��@                           @j���@0           p�@������������������������       ��Cv֯@�           8�@������������������������       ��ꈨO�@�            pp@                           @�)�L-�@�            �t@                            �?_TJ=�@^            �a@                            �?w��C>�@8            �T@������������������������       �.���^@            �D@������������������������       �ig��"�@             E@                           �?�v=�E	@&             M@������������������������       �N�M�t�@             9@������������������������       ��n�� �@            �@@                           @� �OA@x            �g@                            �?@W(��I@^            �a@������������������������       ��<)r6@,            �O@������������������������       �Ҋ���@2             T@                          �=@�$9R� @            �F@������������������������       �EA��W�?             *@������������������������       ��})@             @@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     @r@     ��@      ?@     �M@     �{@     @T@     ��@     `l@     ��@     �x@      =@      0@      p@     �@      <@     �H@     �x@     �P@     ��@      i@     ��@     �s@      :@      @     �S@      i@      @      ,@     �\@      0@     ~@      S@     `t@     @`@      @              <@      L@                      @@      �?     @n@      4@     �`@      E@       @              7@     �F@                      =@      �?     `i@      $@     @U@      ?@       @              @      &@                      @             �C@      $@      I@      &@              @     �I@      b@      @      ,@     �T@      .@     �m@      L@     �g@      V@      @      @      *@      N@       @      @      6@      �?     �X@      .@      U@      @@                      C@      U@      @      &@      N@      ,@     �a@     �D@     �Z@      L@      @      (@     `f@     �s@      7@     �A@     `q@      I@     `}@     @_@     �{@     @g@      5@      (@     �a@      g@      0@      :@      i@      A@     �g@     �Y@     `j@     @_@      *@      @      1@     �L@      @      $@      Q@      @     @Q@      6@     @P@      C@      @      "@      _@     �_@      *@      0@     �`@      <@     �^@     @T@     @b@     �U@      "@              C@     @`@      @      "@     �S@      0@     pq@      6@     �l@     �N@       @              5@     �Y@       @       @      I@      (@      j@      *@     `d@     �A@                      1@      ;@      @      �?      <@      @     �Q@      "@     �P@      :@       @      @      A@     �H@      @      $@     �I@      .@      9@      :@      ?@     �S@      @       @       @      3@      @       @      .@      @      (@      *@      (@     �E@       @              �?      $@              @      @      @      "@       @      @     �@@       @                      "@              �?      @      �?      @       @      @      $@       @              �?      �?              @      �?      @       @      @       @      7@               @      @      "@      @      @      "@              @      @      @      $@               @      �?      @       @      @      @              �?              @      @                      @      @      �?      �?      @               @      @      @      @               @      :@      >@               @      B@      &@      *@      *@      3@     �A@      �?       @      5@      4@               @      8@      &@      @      *@      *@      >@      �?      �?       @      @                      @      @       @      "@      "@      2@      �?      �?      *@      0@               @      4@      @      @      @      @      (@                      @      $@                      (@              @              @      @                              @                      @               @               @                              @      @                      "@              @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�;k�`6@�	           ��@       	                    �?'���		@�           �@                           �?l_�J��@/           0}@                          �6@�����@q            �f@������������������������       ��W��*d@G            @[@������������������������       �D�٢��@*            �Q@                          �3@b�%W�L@�            �q@������������������������       �t5e7n@;            �T@������������������������       ���0�I@�            �i@
                          �2@�qS�u	@�           ȑ@                            �?�O�o��@�            �k@������������������������       �n�5�ko@$             O@������������������������       ���>A��@g            �c@                           �?�D��B�	@6           ��@������������������������       ��H�@�            @u@������������������������       ��AZ�
@q           �@                           �?�n!��@�           �@                            �?5�{�v�@�           (�@                          �8@a�Ow��?r            �f@������������������������       ���ɷ���?f            �c@������������������������       ����D3l@             5@                          �8@x=��@f           ��@������������������������       �k,��e@,           p}@������������������������       �
#v�+@:            �V@                           @N����@�           |�@                            @�SK='�@           �{@������������������������       �.�`Z�@�            Pr@������������������������       ��Dy}��@Z            `b@                           @l���F!@�           ��@������������������������       ������@�           �@������������������������       ��w:���@            �E@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �t@     `�@      A@      M@     �{@     @Q@     Ў@     �i@     �@     �v@      ;@      *@     @h@     �l@      8@      >@     �n@      A@     �k@     `a@     @p@     `h@      4@      @      L@     �R@      �?      @     �M@      @     �Y@      ,@     �X@      G@      @      @      5@      7@                      5@             �J@       @      E@      *@      �?              @      2@                      @              C@       @      @@      @              @      .@      @                      ,@              .@              $@      @      �?             �A@      J@      �?      @      C@      @     �H@      (@      L@     �@@       @               @       @              �?      @       @      ;@       @      (@      .@                      ;@      F@      �?      @      ?@      �?      6@      $@      F@      2@       @      "@     @a@     `c@      7@      8@      g@      ?@      ^@     @_@     @d@     �b@      1@       @      5@      :@      @      @     �C@              E@      <@     �A@      4@      �?              @      @                       @              (@      (@      1@              �?       @      0@      3@      @      @      ?@              >@      0@      2@      4@              @     @]@      `@      3@      5@     @b@      ?@     �S@     @X@     �_@      `@      0@              4@      J@       @       @     �P@      @      C@     �B@     �L@     �I@      @      @     @X@     @S@      1@      *@      T@      9@      D@      N@     �Q@     �S@      *@             �`@     `t@      $@      <@     �h@     �A@     ��@     �P@     �@     �d@      @              @@      W@                     �D@      $@     @t@       @      i@      ?@       @              �?      2@                      ,@      @      X@             �D@      @      �?              �?      .@                      *@             �V@             �A@      @                              @                      �?      @      @              @       @      �?              ?@     �R@                      ;@      @     �l@       @      d@      9@      �?              =@      Q@                      8@      @     `h@      @     �`@      ,@      �?               @      @                      @      @     �@@      @      :@      &@                     �Y@     @m@      $@      <@     `c@      9@     �{@     �M@     @w@      a@      @             �A@      U@      �?      $@      L@      (@     �V@      A@      R@     �F@      �?              5@     �F@               @     �F@      &@     �J@      ;@     �K@      ;@      �?              ,@     �C@      �?       @      &@      �?     �B@      @      1@      2@                      Q@     �b@      "@      2@     �X@      *@     �u@      9@     �r@     �V@      @             �M@     �b@      "@      ,@     @X@       @     �u@      4@      r@      V@      @              "@       @              @       @      @      @      @      $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJZo�~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�b@�O@�	           ��@       	                    �?
��bt@           ��@                            �?)�?�Z�@�           ؄@                            �?�D���@�            �w@������������������������       ��r�l'@d            `d@������������������������       �\/�U@�             k@                          �5@Η�� �@�             r@������������������������       �~{g��@r            �f@������������������������       �+�Ak8"@G            �Z@
                           @t�@n           X�@                            �?�JxiM@�             u@������������������������       ���}9�h@            �i@������������������������       �O@m���@U             `@                          �2@���A� @�            `o@������������������������       ��x} 1B�?>            @X@������������������������       ��?|�@\            @c@                           @���H@�           Ƥ@                          �4@Cƛu�@�           �@                           @��xt@�           T�@������������������������       �q�!/�v@J           �@������������������������       �~��w@V           ��@                           �?O�����@/           ��@������������������������       �P�&���@H             [@������������������������       ��πws�@�           0�@                           @��&Q	@�            `u@                          �3@�
MM�	@s            @h@������������������������       ��l|��@            �A@������������������������       �H!{S�;	@\            �c@                            �?�	���@^            �b@������������������������       ���*�@3             S@������������������������       �[6�q��@+             R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     �s@     ��@      =@     �N@     pz@     @R@     ��@     �h@      �@     �v@      ?@       @     @V@     �f@       @      $@     �X@      $@     �|@     �A@     �p@     �V@      @       @     �C@      X@      �?      "@      L@       @     @p@      6@      _@     �H@      �?       @      5@      L@      �?      "@      >@      @     @c@      $@      M@      A@      �?       @      @      5@              @      &@       @     @S@      @      <@      "@                      1@     �A@      �?      @      3@      �?     @S@      @      >@      9@      �?              2@      D@                      :@      @     �Z@      (@     �P@      .@                      &@      0@                      ,@      @     �T@      "@     �B@      @                      @      8@                      (@              7@      @      =@       @                      I@     �U@      �?      �?     �E@       @      i@      *@     `b@     �D@      @              E@      H@              �?     �B@              T@      &@     @U@      >@       @              =@      9@              �?      *@              E@      @      R@      2@       @              *@      7@                      8@              C@      @      *@      (@                       @      C@      �?              @       @      ^@       @      O@      &@      �?              �?      @                                     @Q@              4@              �?              @      @@      �?              @       @     �I@       @      E@      &@              9@     �l@     �x@      ;@     �I@     @t@     �O@     P�@      d@     ��@      q@      ;@      1@      h@      u@      8@      I@     @q@     �J@     �~@     �`@     �~@     �m@      ,@       @      Q@     `b@      $@      .@     �Z@      $@     0s@      L@     �l@     �T@      @       @     �B@      O@      "@       @     �S@      @     �Z@      G@     �U@     �L@      @              ?@     @U@      �?      @      <@      @      i@      $@      b@      9@              "@     @_@     �g@      ,@     �A@      e@     �E@     �g@     @S@     p@     @c@      $@      @      ,@      (@               @      4@       @      "@      "@      7@      @      �?      @     �[@     `f@      ,@      ;@     �b@     �D@     `f@      Q@     @m@     �b@      "@       @     �B@      K@      @      �?      H@      $@     �M@      <@     �F@      B@      *@       @      4@      B@              �?      =@      "@      5@      7@      *@      8@      $@      �?       @      @                      "@       @       @      �?      @      @      @      @      2@      @@              �?      4@      @      3@      6@      @      4@      @              1@      2@      @              3@      �?      C@      @      @@      (@      @              @      (@      �?              @      �?      6@      @      4@       @                      *@      @       @              ,@              0@       @      (@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ9�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�F*m@�	           ��@       	                    �?�V�i�@k            �@                           �?�,�/9g@�           h�@                           �?J�f�9@�            0q@������������������������       �K�.�F�@U            ``@������������������������       �`�J�R	@\             b@                            �?��� � @3           �}@������������������������       �rM?	�@^             a@������������������������       �� ��@�             u@
                           @���l.�@�           L�@                           �?��׶�H@�           H�@������������������������       ����v@�             p@������������������������       ��۪K�@�            pv@                           @x�JK��@           P�@������������������������       �b���� @E           �@������������������������       ��n���@�            �r@                           �?��90�@U           $�@                           �?��+p�@            �{@                            �?��?�@�            @l@������������������������       �)��>�@S            �`@������������������������       ��)��y@D            �V@                          �=@l%>��@�            `k@������������������������       �J���t�@x            �h@������������������������       ��J��^O@             6@                           @�I�0�	@5           0�@                          �9@jf`wE�	@           @�@������������������������       �Z�W5R;	@           @|@������������������������       �MY>.��	@�            @x@                          �8@��`�|)@*           @|@������������������������       �:�0�@�            @o@������������������������       ���LC@�            @i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     Pr@     ��@      ;@     �K@     �|@     �X@     ��@     �j@     p�@     �v@     �A@      &@     �]@     Pu@      "@      <@     �j@      B@     ��@      T@     �~@     @e@      1@      &@      O@      \@       @      .@     �]@      1@     �`@     �I@     `a@      T@       @      @      <@      I@       @      @      H@      @      K@      7@      C@      .@      @              @      :@      �?       @      <@       @     �@@      @      5@      @              @      6@      8@      �?       @      4@      @      5@      0@      1@      $@      @      @      A@      O@              &@     �Q@      (@      T@      <@     @Y@     @P@      @              "@      .@              �?      8@              8@      @      D@      .@       @      @      9@     �G@              $@      G@      (@      L@      6@     �N@      I@      @             �L@     �l@      @      *@     �W@      3@     p�@      =@     v@     �V@      "@             �@@     �[@       @      @      L@      1@     �h@      4@     �`@      C@      @              *@     �B@               @     �@@      .@     @T@      $@     �E@      4@      @              4@     @R@       @       @      7@       @     �]@      $@     �V@      2@                      8@     �]@      @      "@     �C@       @     pt@      "@     `k@      J@      @              .@     �O@       @      @      2@             �l@      @      b@      >@                      "@      L@      @      @      5@       @     �X@      @     �R@      6@      @      @     �e@     �o@      2@      ;@     `n@      O@      t@     �`@      r@      h@      2@             �C@      Q@      �?      @     �K@      @     �[@      .@     @W@      H@      @              <@      E@              @      A@      �?      7@      "@     �E@      C@      @              4@      6@              �?      .@      �?      $@      @      >@      <@      @               @      4@              @      3@              *@      @      *@      $@                      &@      :@      �?              5@      @     �U@      @      I@      $@      �?              &@      9@      �?              1@      @     �T@      @      G@      @                              �?                      @      �?      @      @      @      @      �?      @     �`@      g@      1@      6@     �g@     �K@     �j@     �]@     �h@      b@      ,@      @     �X@     ``@      (@      1@      _@     �G@     �S@     �Z@     �Z@     �Y@      *@       @      K@     �T@      "@      (@     �Q@      *@      F@     �I@     @P@      E@      @      @     �F@      H@      @      @     �J@      A@      A@     �K@     �D@      N@      @              B@     �J@      @      @      P@       @     �`@      *@     �V@      E@      �?              2@      =@       @      �?      ?@      @     �X@       @      E@      4@      �?              2@      8@      @      @     �@@       @      B@      &@     �H@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO�ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��˗%M@�	           ��@       	                    �?�E���@           ��@                          �6@��ss`@�           h�@                           �?�n�#[@           �z@������������������������       ���م@F            �[@������������������������       �6��Cw @�            �s@                            �?#����Y@~            @h@������������������������       ������@!            �G@������������������������       ����os0@]            `b@
                          �5@��<n�F@�           ��@                           @G*N���@�            �u@������������������������       �FE���@~            @i@������������������������       ��'ɕL�?g            @b@                            @����\@�            �n@������������������������       ��H�@t            @f@������������������������       ��q	p�`@'             Q@                          �5@�~�o64@�           �@                           �?YF��\�@�           ��@                           �?���Rw	@Q           8�@������������������������       ��\���\@�            @i@������������������������       �p�B2�	@�            �s@                           �?���ذ�@9           Ќ@������������������������       ������@           @z@������������������������       ��q�-�@5           `@                           @�Q�RC3	@            ��@                           @ւd��	@           ��@������������������������       �2�*�ж	@�            �@������������������������       �c?PŜ@M             ]@                           @e�R|��@           {@������������������������       �V��F@�            �r@������������������������       ����^�
@]             a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     t@     ��@     �A@     �O@     `z@     �T@     ��@     �h@     8�@     �v@      9@      �?     @Q@     @e@       @      ,@      Y@      &@      {@      H@     �q@     @S@      @      �?      <@      T@      �?      *@     �N@      "@     �n@      6@     �^@      B@                      .@     �K@              @      @@      @     `i@      *@     @T@      1@                       @      &@              @      ,@       @      A@      $@      3@       @                      @      F@              @      2@       @      e@      @      O@      "@              �?      *@      9@      �?      @      =@      @      F@      "@      E@      3@              �?      @      @               @      @      @      *@      �?      @      @                      $@      2@      �?      @      7@              ?@       @      C@      ,@                     �D@     �V@      �?      �?     �C@       @     `g@      :@     `d@     �D@      @              6@      L@                      (@              b@      @     @V@      3@                      ,@      B@                      &@              N@       @     �O@      0@                       @      4@                      �?              U@      @      :@      @                      3@      A@      �?      �?      ;@       @     �E@      4@     �R@      6@      @              *@      4@      �?      �?      6@       @      :@       @     �P@      .@      @              @      ,@                      @              1@      (@      @      @              2@     �o@     �x@     �@@     �H@      t@     �Q@      �@     �b@     H�@     �q@      6@      "@     @Y@      k@      ,@      6@     �b@      ;@     �x@     �J@     @t@      ^@      $@      "@     �M@     �S@       @      "@     @V@      3@      O@     �@@     �S@     @P@      "@      �?      (@      A@              @     �@@      @      A@      "@     �A@     �@@               @     �G@      F@       @      @      L@      ,@      <@      8@      F@      @@      "@              E@     @a@      @      *@      N@       @     �t@      4@     �n@     �K@      �?              5@     �M@      @       @     �C@      @      a@      @     �\@      ;@      �?              5@     �S@      �?      @      5@      @     �h@      ,@     ``@      <@              "@     �b@     �f@      3@      ;@     �e@      F@      g@      X@     �h@     �d@      (@      "@     @[@     �`@      .@      4@      ^@     �D@      T@     �R@     �X@     �[@      (@      @     �X@     @\@      *@      4@     �[@      B@     �P@     �I@     @V@     @W@      &@      @      $@      6@       @              $@      @      *@      7@      "@      2@      �?              E@      G@      @      @     �J@      @      Z@      6@     �X@     �J@                      9@      ?@       @      @      C@              V@      &@      Q@      ?@                      1@      .@       @      @      .@      @      0@      &@      ?@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�# hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @� �}0@�	           ��@       	                   �7@v�����@|           \�@                           �?v��8�@�           ��@                           �?n0"��<@�           ��@������������������������       �0��ž�@�             t@������������������������       �� �a��@�           ��@                            @9�w�:@�            Px@������������������������       ���s�%�@�            Pr@������������������������       ��?�$�@E             X@
                           �?r�(>�	@�           ��@                          �<@z�>��@�            �l@������������������������       ��Y�;^�@c            �d@������������������������       �]l�9�@(            @P@                           �?<�A���	@p           X�@������������������������       �L����C@u            �g@������������������������       ��^V�	@�            �x@                            @�;�M�@4           l�@                           �?ϗ�t/�@�           ��@                            �?����$@�           �@������������������������       �����6�@&           �|@������������������������       ��-s)V@�            �n@                           @yi"A��@�           @�@������������������������       ��zw���@�            �s@������������������������       ��ܙ��@�             w@                           �?���m� @�            s@                           �?�q�.{�??            �\@������������������������       �[���
�?)             S@������������������������       ��h��?��?            �C@                           @���W@t            �g@������������������������       ���%�X��?>            @Z@������������������������       ������@6            @U@�t�b�~     h�h5h8K ��h:��R�(KKKK��h��B�        *@      t@     ؁@      =@      I@     P|@     @W@     `�@     �j@     `�@     �t@      8@      (@     `n@     0t@      7@     �B@     �s@      S@     �v@     �f@     @x@      n@      3@      @     �`@     �l@      @      8@     �h@      B@     p@     �Y@     �q@      ]@       @      @     @\@      e@      @      3@     �b@      ;@     �b@     �S@     �i@     �W@      @             �D@      K@              �?     �@@      @     �O@      1@     �T@      :@              @      R@     �\@      @      2@     �\@      7@     @U@     �N@     @^@      Q@      @              6@      O@       @      @     �I@      "@     @[@      8@     �T@      6@      �?              5@      G@       @       @      D@      @      S@      1@     �Q@      *@      �?              �?      0@              @      &@      @     �@@      @      (@      "@              @      [@     @W@      1@      *@     �]@      D@     �Z@     �S@     �Y@      _@      &@      @      ;@      <@       @      �?      >@      @     �C@      ,@      D@     �A@      @      @      ,@      2@      �?              ;@      �?     �A@      @      >@      7@      @              *@      $@      �?      �?      @      @      @      @      $@      (@               @     @T@     @P@      .@      (@      V@     �A@      Q@      P@      O@     @V@      @      �?      @@      3@               @      @@      @      7@      5@      4@      <@              �?     �H@      G@      .@      @      L@      ?@     �F@     �E@      E@     �N@      @      �?     @S@      o@      @      *@      a@      1@      �@      A@     �z@     �V@      @      �?      Q@      m@      @      (@     �Y@      .@     �~@      @@     �u@     @R@      @      �?     �B@     @_@       @      $@     �N@      @     0p@      *@      c@      C@       @              5@      T@      �?       @      D@      @     `e@      @      Z@      8@      �?      �?      0@     �F@      �?       @      5@              V@      @      H@      ,@      �?              ?@     �Z@       @       @      E@      "@     �l@      3@     �h@     �A@      @               @      K@      �?       @      .@       @     @[@      .@     �U@      (@      �?              7@     �J@      �?              ;@      �?     �^@      @      \@      7@       @              "@      0@       @      �?     �@@       @     �b@       @     @R@      1@                      @      �?                      @             @U@              3@      @                      @                              @             �I@              .@      @                              �?                                      A@              @                              @      .@       @      �?      >@       @     @P@       @      K@      ,@                              @                      3@      �?     �E@      �?      A@      �?                      @      "@       @      �?      &@      �?      6@      �?      4@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@Ȉ��x@o	           ��@       	                    �?��t@8           �@                           �?�Gä�J@�           ��@                           �?6�,�f@�            `p@������������������������       �r1�	-@M             _@������������������������       ����U�@R            @a@                            �?}�y5^	@+            }@������������������������       �!�}�@X             b@������������������������       �fr���?	@�            �s@
                           @Y��M@n           ��@                           �?�s�}@y           �@������������������������       �wWԧ�@�            @m@������������������������       �����;2@�            py@                           @.��yMr@�           `�@������������������������       �ڪ��> @?            �@������������������������       �.�1�	@�            �r@                            �?3�(qhX@7           �@                          �6@��	@�@%           ��@                           �?�c�(5!@^            �b@������������������������       �S���Gi@(            �O@������������������������       �:��5F�@6            �U@                           �?j��i��@�           �@������������������������       ����ƻ�	@�            pv@������������������������       ����>�@�            �w@                          �<@�Ơr�@           ��@                           @9��m�@@�           ��@������������������������       �6�J�@�           0�@������������������������       ������@-             S@                            @�ӢH#	@`            �c@������������������������       �����;x@             A@������������������������       �6~(�	@L             _@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     `r@     h�@      :@     �H@     �|@     @P@     T�@     �i@     �@     @v@      >@      "@     �^@     �r@      @      7@     �j@      <@      �@     �T@     0~@     `d@      .@      "@     �O@      Y@      @      (@      Y@      ,@      b@      H@     `a@      U@      $@              1@     �G@      �?       @      5@      �?     @T@      ,@     �K@      5@       @              @      2@      �?              .@      �?      D@       @      3@      *@       @              $@      =@               @      @             �D@      @      B@       @              "@      G@     �J@       @      $@     �S@      *@     �O@      A@      U@     �O@       @              *@      2@              �?      4@      @      :@      "@      B@      *@      @      "@     �@@     �A@       @      "@     �M@      $@     �B@      9@      H@      I@       @              N@     �h@      @      &@      \@      ,@     ��@     �A@     �u@     �S@      @              B@     @Z@      @      @      L@      ,@     �k@      9@      a@      D@       @              2@      A@                      @       @     �W@       @     @P@      (@                      2@     �Q@      @      @     �H@      (@     �_@      7@     �Q@      <@       @              8@      W@      �?      @      L@             @w@      $@      j@     �C@      @              &@     �M@      �?      @      :@             @p@      @     �_@      6@                      *@     �@@               @      >@              \@      @     @T@      1@      @      $@     `e@     @p@      3@      :@     `o@     �B@     Ps@     �^@      t@      h@      .@      @     �U@      ^@      @      0@     �^@      ;@      d@     �P@     �c@     �Z@      &@       @      3@      >@       @      @      .@      @     �D@      @      3@      $@                      @      &@              �?      &@              :@              @       @               @      (@      3@       @      @      @      @      .@      @      ,@       @              @     �P@     �V@      @      (@      [@      8@     �]@      O@     `a@     @X@      &@      @      B@     �D@      @      "@      O@      &@     �B@      D@      J@     �J@      $@              ?@     �H@              @      G@      *@     �T@      6@     �U@      F@      �?      @     @U@     �a@      ,@      $@      `@      $@     �b@     �L@     @d@     �U@      @       @     @Q@     �\@       @      @     @X@      @     �`@      E@     @b@     �O@      @       @      N@      X@      @      @     �U@      @     @]@      A@     �a@      M@      @              "@      2@      @              &@       @      1@       @      @      @              �?      0@      :@      @      @      ?@      @      .@      .@      0@      7@                      @      @                      .@       @      @              �?       @              �?      &@      7@      @      @      0@       @      "@      .@      .@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��PhhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�D512t@�	           ��@       	                    �?![D�|�@�           N�@                           �?���.�1	@           (�@                           �?��4�ڎ@:           �}@������������������������       �����r@�            �l@������������������������       �����F/@�             o@                           �?JC���	@�           ��@������������������������       �,��#�I@           �y@������������������������       �)웞O
@�           ��@
                           �?� ��@�           �@                          �2@�Yb�@r            �f@������������������������       ��.[��h @&             P@������������������������       ��\����@L            �]@                           �?' ��S@           pz@������������������������       ����p�@f            �d@������������������������       ����2@�            p@                          �7@����$@!           ��@                           @rDt��@           (�@                           �?���?�A@3           ��@������������������������       ��!|�g@-            ~@������������������������       ��Y�]<� @           �z@                            �?�c���@�            �w@������������������������       �V�G|��@1             U@������������������������       �E��0�9@�            `r@                            �?oΔ^��@           �y@                           @|�-j�@�            @j@������������������������       �ET�<e@U            �`@������������������������       �C��@-            �S@                           @v|]���@�            �h@������������������������       � �؊@?            �X@������������������������       �{�R�C@B            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �r@     h�@      @@     �O@     P}@     �V@     ��@     �j@     ��@     @v@      9@      7@     @i@     Pu@      7@     �E@      t@     �Q@     �v@     �f@      w@     �o@      4@      7@     @c@     �n@      6@      <@     `o@      H@     �k@     �`@     pp@     `i@      3@      �?     �B@      S@              @     @P@      @      Y@      9@     �Z@     �L@       @      �?      2@      @@              @      <@      @     �K@      .@     �C@      ?@       @              3@      F@              �?     �B@             �F@      $@     �P@      :@              6@     @]@     @e@      6@      7@     @g@      F@     @^@     �Z@     �c@     @b@      1@       @     �@@     �Q@      @       @      T@      @      O@      ?@     �K@     �I@      @      4@      U@     �X@      1@      .@     �Z@     �C@     �M@      S@     �Y@     �W@      (@              H@     �W@      �?      .@     �Q@      7@      b@      I@     �Z@      I@      �?              4@      5@              �?      .@       @     �Q@      @     �C@      @                       @       @                      @              =@              1@      @                      2@      *@              �?      $@       @      E@      @      6@      @                      <@     �R@      �?      ,@      L@      5@     @R@     �E@      Q@      F@      �?              "@      <@      �?       @      <@       @      9@      $@      ?@      7@      �?              3@      G@              (@      <@      *@      H@     �@@     �B@      5@               @     @Y@      k@      "@      4@     `b@      3@     ��@      ?@     @x@     �Y@      @             @Q@     �e@      @      (@     �V@      *@     ��@      (@     �q@     �P@      @             �D@     �\@       @             �H@      @     @{@       @      j@     �F@      �?              <@     �G@                     �D@      @     `m@      @      Y@      7@      �?              *@     �P@       @               @      @      i@      @     @[@      6@                      <@     �N@      @      (@     �D@      @     @_@      @     @R@      6@       @              @      "@       @      �?      @       @      F@              (@      @                      9@      J@       @      &@      A@      @     @T@      @     �N@      2@       @       @      @@     �D@      @       @     �L@      @      X@      3@     �Z@      B@       @              8@      9@              @      9@      @     �G@      "@     �H@      4@                      $@      6@              @      *@      @      D@      @      6@      &@                      ,@      @                      (@      @      @      @      ;@      "@               @       @      0@      @      @      @@             �H@      $@     �L@      0@       @       @      @      @              �?      7@              7@      @     �@@      @       @              @      &@      @       @      "@              :@      @      8@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�c1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @T;V�@�	           ��@       	                    �?�L:��	@]           >�@                          �;@9�UzJ�@�           H�@                           �?t#��9�@g           ��@������������������������       ���\��,@           �y@������������������������       �@���@f             c@                           �?�4έS@5            �T@������������������������       ����7��@,            �P@������������������������       ��u�B�+@	             .@
                           �?:�7S�	@�           X�@                          �2@UB�\]�	@�           `�@������������������������       ���b��9@            `j@������������������������       ���ަ�>
@B           (�@                           �?�wɵ��@            �w@������������������������       �ϲ���I@            �@@������������������������       �_�	>~@�            �u@                          �5@�O�Z)*@9           ��@                           �?a�B�qx@�           D�@                          �0@n&�'{8�?�            x@������������������������       �@�Y�?            �J@������������������������       ��y7����?�            �t@                           @c9���@�           ��@������������������������       �l=x�(@}           @�@������������������������       �{�,�~@)             R@                           @�`WF@�           Ȅ@                           �?�� ��@�           8�@������������������������       ��R�;O@�            �s@������������������������       �d>�;��@�            �t@������������������������       ��Yk�M@             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        7@     �s@     (�@      @@     �K@     �y@     �U@     x�@      n@     ��@      w@      =@      7@     `l@     ps@      5@      F@     �r@      O@      w@     �i@      x@     `m@      :@      �?     @R@     @U@              (@     �Q@      @      c@     �C@     �c@      I@      @             �P@     @R@               @     �I@      @     �b@     �@@      b@      B@      �?              L@      N@              @     �B@       @     @Y@      @@     @W@      ;@      �?              $@      *@               @      ,@       @      I@      �?     �I@      "@              �?      @      (@              @      3@       @       @      @      (@      ,@      @      �?      @      (@              @      (@       @       @      @      $@      *@                      �?                              @                      �?       @      �?      @      6@     @c@     @l@      5@      @@     �l@      L@     �j@     �d@     �l@      g@      6@      6@     �\@     @c@      4@      ;@     �f@     �D@     `b@     @`@      e@     �b@      5@      @      0@     �B@              @     �A@              A@      1@     �C@      :@      �?      3@     �X@     @]@      4@      8@     `b@     �D@     @\@     @\@      `@     �^@      4@             �C@      R@      �?      @      H@      .@      Q@     �B@      N@      B@      �?              @      @              @      @      �?      �?      "@      @      @                      A@     @Q@      �?       @     �F@      ,@     �P@      <@      L@      @@      �?              W@     �m@      &@      &@     �\@      9@     ��@     �A@     @{@     �`@      @              E@      c@      �?      @     �E@      .@     Pz@      (@     �q@     @P@       @              &@      L@              �?      (@      �?     `i@      @      U@      *@                              *@                       @              =@              @      @                      &@     �E@              �?      $@      �?     �e@      @      T@       @                      ?@     @X@      �?      @      ?@      ,@     @k@       @     �h@      J@       @              9@     �V@      �?      @      <@      "@     @h@      @      g@      C@       @              @      @               @      @      @      8@      �?      &@      ,@                      I@     @U@      $@      @      R@      $@     @g@      7@     �c@      Q@      �?              F@      U@      @      @     �P@      "@     @g@      5@     �c@      Q@      �?             �@@      F@      �?      @      >@      @      Y@      @      Q@      9@      �?              &@      D@      @      �?     �B@      @     �U@      0@      V@     �E@                      @      �?      @              @      �?               @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�+�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @gZ��p@�	           ��@       	                     @T^�7z�@w           ��@                           �?�(�,�@x           ��@                          �<@N:��o	@[           ��@������������������������       ��6%��@           ��@������������������������       �T{�5�@N            @`@                           �?��v�N@           �}@������������������������       ��<k��@R            `a@������������������������       �����@�            �t@
                          �1@NO:��	@�           ��@                           �?��O@G            �\@������������������������       �NZk@6             V@������������������������       ����|���?             :@                           �?����L	@�            �@������������������������       �����	@�             q@������������������������       ���+��k@            y@                          �7@a�̅@;           $�@                           �?�H�¿�@5           $�@                           �?+�!uD @%           �z@������������������������       ���}e��?�            �n@������������������������       �ʕ��� @{             g@                           @�|P�ų@           �@������������������������       �$w��@            �j@������������������������       �������@�           0�@                           �?45	[ �@            x@                            @ߞ[�?�@}            @g@������������������������       �E�ƣL�@l            @d@������������������������       ��I
Ւ @             8@                           @F��D@�            �h@������������������������       ����K�@=            �U@������������������������       ����ǉ@L             \@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     0q@     �@      A@      L@     �~@     @W@     ��@     `m@     ��@      v@      9@      2@     �g@     �t@      8@      I@     �u@     �R@     �v@     `h@     pw@     �n@      2@       @     �\@     �i@      $@     �A@      n@      H@     `o@     �a@     �l@     �c@      &@       @      U@      a@      "@      9@     �f@      @@     �a@     �W@     �`@     @_@      $@      @      R@     �_@      "@      8@     �d@      5@      a@      T@     �\@      V@      "@      �?      (@      $@              �?      1@      &@      @      ,@      3@     �B@      �?              >@     @Q@      �?      $@      M@      0@      [@     �H@     �X@     �@@      �?               @      1@              �?      *@      @      K@      @     �@@      @                      6@      J@      �?      "@     �F@      *@      K@     �E@     @P@      =@      �?      $@      S@      `@      ,@      .@     �[@      ;@     @\@      J@      b@      V@      @              &@      0@      �?      �?      (@              A@       @      1@      ,@                      $@      "@      �?      �?      (@              7@      @      *@      ,@                      �?      @                                      &@      @      @                      $@     @P@     @\@      *@      ,@     �X@      ;@     �S@      F@     �_@     �R@      @      @     �A@     �E@      $@      $@      F@      .@      <@      @      E@      ?@       @      @      >@     �Q@      @      @     �K@      (@     �I@      C@     @U@     �E@      @       @     @U@     �j@      $@      @      b@      2@     H�@      D@     pz@      [@      @              K@     �e@      @      @      W@      *@     ��@      1@     `s@      R@      @              .@      H@       @       @      4@       @      m@       @     @V@      "@      �?              @      6@               @      .@       @     �a@       @     �G@      @                       @      :@       @              @              W@      @      E@       @      �?             �C@     @_@      @      �?      R@      &@     `s@      "@     �k@     �O@      @              &@      B@      �?              0@      &@     @Q@      @      F@      2@      @              <@     @V@      @      �?      L@              n@      @      f@     �F@      �?       @      ?@      D@      @      @      J@      @     �R@      7@     @\@      B@      �?       @      4@      9@              @      4@              >@      $@      P@      &@      �?       @      4@      6@              @      3@              3@      "@      M@      "@      �?                      @                      �?              &@      �?      @       @                      &@      .@      @              @@      @     �F@      *@     �H@      9@                       @      $@       @              $@      @      5@      "@      1@      $@                      "@      @      �?              6@              8@      @      @@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ/�N hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?r��P@�	           ��@       	                    �?��7'�@	           ,�@                          �<@�g��@6           �}@                           �?�B���v@           �y@������������������������       �w� T�4@a             c@������������������������       �%`��s�@�            0p@                          @@@s���S�@*            @P@������������������������       ����s�`@"             J@������������������������       �V@���@             *@
                           �?I��b@�           x�@                          �;@ �n���@           �y@������������������������       �����2@�            px@������������������������       �;�5�;@             1@                            @f��p@�            pu@������������������������       � ,U{��@�            �q@������������������������       ���)�>��?%             M@                          �5@j���$@�           ��@                           �?��?;bc@�           �@                          �4@G�0�`8@4           �}@������������������������       �m�1��@�            �w@������������������������       ��j�3�@<            �W@                          �3@:\�W�t@Q           `�@������������������������       ��Ku�S@�           `�@������������������������       ����l�@�             t@                           @�pZW	@           ��@                          �;@�΢���	@            �@������������������������       ��>>!�B	@v           ��@������������������������       ���L�
@�            �n@                           �?s��p�@           @{@������������������������       � ���,2@             5@������������������������       ��`'LP�@           �y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@      s@     `�@      =@     �I@     0}@     @S@     �@     �m@     ȉ@     Pv@      5@             @V@     �d@       @      .@     �[@      @     �y@     �G@     �r@     @T@      @              J@     �P@      �?      $@     �N@       @     @V@      :@     @[@     �L@       @              G@     �M@      �?      @      J@       @     �U@      5@     �Y@      @@       @              *@      1@                      1@              D@      �?     �J@      $@      �?             �@@      E@      �?      @     �A@       @     �G@      4@     �H@      6@      �?              @       @              @      "@               @      @      @      9@                      @      @                      @               @      @      @      9@                       @      �?              @      @                              @                             �B@     @X@      �?      @     �H@      @      t@      5@      h@      8@       @              1@     �G@              @     �A@       @     �g@      "@     @V@      *@                      ,@      E@              @     �A@             �g@      @      V@      &@                      @      @                               @       @       @      �?       @                      4@      I@      �?              ,@      �?      `@      (@     �Y@      &@       @              2@     �H@      �?              (@      �?      X@       @     �U@      &@       @               @      �?                       @             �@@      @      0@                      6@      k@     �x@      ;@      B@     Pv@      R@     P�@      h@     `�@     @q@      1@      @     @U@     �i@      $@      ,@     �b@      ;@      w@     �Q@     pu@      a@       @      @      H@     @Q@       @      @      T@      .@     �L@     �B@     @U@     �Q@      �?      �?      F@      E@       @       @     �P@      $@     �H@      @@     @Q@     �N@      �?      @      @      ;@              @      ,@      @       @      @      0@      "@                     �B@     �`@       @      "@     �Q@      (@     ps@     �@@      p@     �P@      �?              6@     �T@      @      @     �A@      @     `m@      7@      e@     �D@                      .@     �J@      @       @     �A@      "@      S@      $@     @V@      9@      �?      1@     �`@     �g@      1@      6@     �i@     �F@     @g@     �^@     �f@     �a@      .@      ,@      X@      `@      *@      3@     �`@      D@      V@      Y@     �W@     �W@      ,@       @      R@     �X@       @      *@      X@      8@     �P@     �S@      R@      J@      "@      (@      8@      =@      @      @     �C@      0@      5@      6@      7@      E@      @      @      B@      N@      @      @      R@      @     �X@      6@     �U@      G@      �?      @       @      �?              �?       @               @      @      @                              A@     �M@      @       @     �Q@      @      X@      1@     @T@      G@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJM�c	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���}y@�	           ��@       	                    @���3`@�           t�@                          �1@��X
��@>           �@                           @���<{�@�             q@������������������������       �M�l�y*@�            0p@������������������������       ���n��S@	             .@                           �?����Jb@�           x�@������������������������       �&U���:@|            �i@������������������������       �kSE��F	@            z@
                          �1@�$�3��@J           ��@                           �?��:��?�             v@������������������������       ��HOϪ @w            `h@������������������������       �s��b��?h            �c@                           @�M��M�@k           ��@������������������������       �W�Y�f@�            �l@������������������������       �uw�@�            Pu@                           @��h�W�@1           X�@                            �?.��(v@�           p�@                           @�j�e@H           ��@������������������������       �g3����@           p{@������������������������       �Y>z���@9            �W@                          �<@�Ü�i@[           �@������������������������       �,�M<�@�           ��@������������������������       ����{	@�            �k@                            �?8]��@�             j@                           �?�oH�@J            �\@������������������������       ��4lX	@             B@������������������������       ������@1            �S@                            @t�6k�@D            @W@������������������������       ��?�s!@             B@������������������������       ��)�>T�@'            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@     X�@      :@     �P@     �y@     �[@     ؏@      k@     �@     �v@     �A@      @      V@     `l@      @      >@     �b@      =@     ��@     @U@     z@      a@      &@      @      M@      _@      @      0@     @Y@      9@     �j@      R@     �f@      U@      $@       @      3@     �@@       @      �?      =@       @     @V@      1@     �L@      7@               @      1@      @@       @      �?      :@             @V@      .@      J@      7@                       @      �?                      @       @               @      @                      @     �C@     �V@      �?      .@      R@      7@     �_@     �K@     �_@     �N@      $@              1@      ?@              �?      4@              J@      *@      L@      0@      �?      @      6@      N@      �?      ,@      J@      7@     �R@      E@     �Q@     �F@      "@              >@     �Y@       @      ,@      H@      @     pz@      *@     @m@      J@      �?              @      D@              @      1@             �g@       @      T@      &@      �?              @      2@              @      *@             �Y@      �?     �C@       @                              6@                      @             @U@      �?     �D@      @      �?              8@     �O@       @      @      ?@      @     `m@      &@     @c@     �D@                      *@     �@@      �?              1@      @     �R@      @     �L@      ;@                      &@      >@      �?      @      ,@      �?      d@      @     @X@      ,@              ,@     �h@     �t@      5@     �B@     �p@     @T@     �w@     ``@      x@      l@      8@      $@     �e@      r@      3@     �B@     `n@      Q@     �u@     �X@     w@     `j@      3@      @      D@      V@      @      @      R@      5@     �Z@      @@     �Y@      G@      $@      @      @@     �Q@      @      @      L@      5@     �U@      ;@     �S@     �F@      $@               @      1@      �?      �?      0@              4@      @      9@      �?              @     �`@      i@      .@      >@     `e@     �G@     @n@     �P@     �p@     �d@      "@      @      [@     �e@      $@      2@     `a@     �A@      l@     �I@      n@     �]@      "@      @      9@      <@      @      (@      @@      (@      2@      0@      9@     �G@              @      :@      D@       @              7@      *@     �@@      @@      1@      *@      @       @      2@      2@      �?              @      $@      1@      9@      $@      "@      �?              $@      @                       @      @      @      @       @                       @       @      *@      �?               @      @      &@      4@       @      "@      �?       @       @      6@      �?              3@      @      0@      @      @      @      @               @      @                      (@      �?      @      �?      @       @      @       @      @      2@      �?              @       @      $@      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJK�@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?.x@K�@�	           ��@       	                    @���?H@�           L�@                           �?�*_@�           ��@                          �6@�$
[j@�             o@������������������������       ��Ot-��@Z            �a@������������������������       �^�����@I             [@                           �?a$�H�<@           �y@������������������������       �φ�[#A@@             Y@������������������������       ������@�            �s@
                           �?/�O�w!@�            �w@                          �5@���j}@v            �g@������������������������       ��`���@O            ``@������������������������       ��{���@'            �L@                           @3g�=U@v             h@������������������������       ���dS]@             H@������������������������       ���4}�g@Y             b@                           @Xc�@&           l�@                          �8@kw���@�           D�@                          �1@�RP��@�           �@������������������������       ��9,MV@t             g@������������������������       �A��@L           H�@                           �?R��8nw	@"           �|@������������������������       � A�ɧ	@�            @w@������������������������       �@ނ6 @7            �V@                           @�|v��@D           ��@                           �?����1!@           �@������������������������       ��b�8r�@5           �~@������������������������       ��ɜ��@�           x�@                            �?�8}&ޏ@@             [@������������������������       ���%�@             C@������������������������       �H�oHBa@'            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     ��@      4@     �H@     �@     @T@     X�@     �i@      �@      u@      :@             �R@      b@      @      &@     �a@      9@     �q@     �P@     �f@     @Y@      &@             �N@     @X@      @      &@     �Z@      4@     @_@     �M@     @Y@      Q@      &@              5@      B@       @      @      D@      @      J@      <@      @@      5@      @              0@      8@              �?      0@      @     �B@      $@      8@       @      �?              @      (@       @      @      8@      @      .@      2@       @      *@      @              D@     �N@      �?      @     �P@      *@     @R@      ?@     @Q@     �G@      @              "@      8@                      $@              3@              >@       @                      ?@     �B@      �?      @      L@      *@      K@      ?@     �C@     �C@      @              *@      H@       @              A@      @     �c@      @     �T@     �@@                      @      5@                      8@       @     �P@      @     �F@      3@                              "@                      1@              J@       @      B@      .@                      @      (@                      @       @      .@       @      "@      @                      @      ;@       @              $@      @     �V@      @     �B@      ,@                      �?      ,@       @              �?              4@       @      @      @                      @      *@                      "@      @     �Q@      �?     �@@      $@              5@     @l@     pz@      .@      C@     �v@      L@     ��@     `a@     H�@     `m@      .@      4@     @d@      n@      (@      :@      p@      E@      m@     �Z@      q@      e@      &@      &@      Z@      e@      @      6@     @g@      5@     �g@     �J@     �k@     �Z@      @      @      @      9@       @      �?      >@              K@      @      E@      ,@               @     @X@     �a@      @      5@     �c@      5@     �`@      G@     @f@      W@      @      "@      M@     @R@      @      @     �Q@      5@     �F@      K@      K@     �O@      @      "@     �F@     �M@      @      @     �O@      1@      ?@      G@     �B@     �H@      @              *@      ,@                      @      @      ,@       @      1@      ,@              �?      P@     �f@      @      (@      [@      ,@     �~@      @@     pu@     �P@      @      �?      H@     �d@      �?      (@     @W@      $@     �|@      <@     �t@      N@      �?              2@     �Q@              �?      :@      @     �k@      &@      ^@      ,@      �?      �?      >@     @W@      �?      &@     �P@      @     �m@      1@      j@      G@                      0@      2@       @              .@      @      :@      @      ,@      @      @              @      $@                              @       @      �?      @      @                      &@       @       @              .@              2@      @       @       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�G6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?E)H�u(@�	           ��@       	                   �8@2@�	@           �@                           �?3��5�Y@�           А@                            @������@           @{@������������������������       �o����@�             r@������������������������       ��(L���@a            �b@                           @��M;L	@�            �@������������������������       �����:�@�           ��@������������������������       ��#��v@            �E@
                           �?�ʿ6U�	@L           p�@                            �?���׃.@S            �^@������������������������       �?���9�@!             J@������������������������       �	���@2            �Q@                           �?���F5�	@�            @y@������������������������       ���>�r�	@\             b@������������������������       �����x	@�            0p@                          �4@ޭ:x�
@�           �@                           �?"�����@            Ԓ@                           @U �j��?           `{@������������������������       �zY���?�            �t@������������������������       �<��!H?@C            �Y@                           @�ߒ'�-@�           ��@������������������������       ��<��@�            �s@������������������������       � $��w@$           @|@                           @^�[�K�@�           H�@                           @m8s��\@2           0~@������������������������       �3M�@�            �s@������������������������       �J΍��@l            �d@                           @nd~\�@~           x�@������������������������       �԰\�N@�            �t@������������������������       �.�|i�T@�            Pr@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     ��@      :@      J@     �|@      T@     H�@     �j@     �@     �v@      =@      (@     �d@      n@      2@      A@      m@     �E@     �n@      a@     p@     �h@      5@      @      ]@      c@      &@      6@      d@      7@     �h@     �Q@     �h@     @[@       @       @      :@     @R@       @       @     @R@       @     �Z@      2@     �T@      D@       @              5@      H@      �?      @     �G@       @      O@      .@     �J@     �@@       @       @      @      9@      �?      @      :@             �F@      @      >@      @              @     �V@      T@      "@      ,@     �U@      5@     �V@     �J@      ]@     @Q@      @      @     @V@     �R@      "@      ,@     �T@      2@      V@      D@     @\@     �N@      @      �?      �?      @                      @      @      @      *@      @       @      �?      @     �I@     �U@      @      (@     @R@      4@     �G@     @P@      M@     �U@      *@              1@      :@              @      3@      �?      *@      @      @      :@       @              @      .@                      @      �?      @       @      @      *@                      &@      &@              @      0@              @      @      �?      *@       @      @      A@     �N@      @       @      K@      3@      A@      M@     �I@     �N@      &@      @      "@      <@      @      @      2@      &@       @      6@      $@      9@       @      @      9@     �@@      �?      @      B@       @      :@      B@     �D@      B@      "@      �?      a@     �r@       @      2@     @l@     �B@     ��@     �S@     ��@      e@       @              P@      c@      @       @     �S@      @     �~@      9@      s@      R@       @              3@      E@               @      ,@             `k@      @      ^@      1@       @              (@      <@                      $@              g@      �?     �U@      *@                      @      ,@               @      @              A@       @      A@      @       @             �F@     �[@      @      @     @P@      @     �p@      6@     @g@     �K@                      7@     �L@      �?      @     �A@       @     @W@      4@     �L@      8@                      6@     �J@      @      @      >@      �?      f@       @      `@      ?@              �?      R@     �b@      @      $@     `b@      A@     �p@     �J@     �p@      X@      @      �?      D@     �J@              @     �R@      9@     @]@      A@     @W@     �C@      @             �@@      B@               @     �G@      .@     �P@      >@      M@      :@      @      �?      @      1@              �?      ;@      $@      I@      @     �A@      *@      �?              @@     �X@      @      @     @R@      "@     �b@      3@     �e@     �L@       @              .@      G@                      B@              X@      @      Y@      ?@                      1@      J@      @      @     �B@      "@      K@      *@     @R@      :@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�aihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�7%�%.@�	           ��@       	                   �5@�<	<�C@	           ē@                           �?ê�j�0@�           ��@                          �3@���	��@�            �n@������������������������       �q�<`Ů@g             d@������������������������       ���->5g@/            @U@                          �3@��)l� @L           ��@������������������������       ����
 @�            �w@������������������������       �.]�S�� @`            �d@
                          �8@���;J@'           �}@                           �?c���H@�            �k@������������������������       �g� :v@?            @Z@������������������������       �� ��@J            �]@                          �<@�K�@�             p@������������������������       ���f�i@d            �d@������������������������       �!����@:             W@                           @*m�ϐ'@�           ��@                            �?��ˇ�O	@�           ȗ@                           �?��ÀJT	@�           ��@������������������������       �C���@�             o@������������������������       ��(䧈�	@X           8�@                           �?4:�	@�           ��@������������������������       ��:��H\	@f           �@������������������������       �U���@{             f@                          �4@����@�           ��@                           �?*(�>�?@o           �@������������������������       �^J�@�            �q@������������������������       �Z "�	D@�            �r@                           @���ځ�@e           �@������������������������       �j��i@2           `}@������������������������       �~���@	@3            @S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     r@     �@     �@@     �H@     P}@     �U@     ��@     �h@      �@     v@      <@              T@      f@      @       @     @[@      (@     P}@     �D@     �q@     �R@      @             �E@     �W@      @      @     �G@      @     �u@      8@     �e@      C@      @              <@      A@      @      @      4@      @     �O@      2@      M@      (@       @              *@      6@                      3@      @     �E@      (@      C@      $@                      .@      (@      @      @      �?              4@      @      4@       @       @              .@      N@              @      ;@      @     �q@      @     @]@      :@       @              (@      B@                      .@              h@      @     �W@      3@       @              @      8@              @      (@      @     @V@      �?      6@      @                     �B@     �T@              �?      O@      @     @_@      1@      \@     �B@      �?              6@      A@                      ?@              Q@      @     �I@      *@      �?              1@      ,@                      5@              1@      @      8@       @      �?              @      4@                      $@             �I@              ;@      @                      .@      H@              �?      ?@      @     �L@      ,@     �N@      8@                      @      =@              �?      3@      @     �D@       @      G@      "@                      "@      3@                      (@              0@      @      .@      .@              4@      j@     �v@      >@     �D@     �v@     �R@     �@     �c@     �@     `q@      7@      3@     �a@     �k@      2@      =@      o@      N@     `j@     �`@     �k@     �h@      1@      @     �T@     @^@      @      6@      [@     �B@     @]@     �P@     �^@     �Y@      @       @      3@     �D@      �?      @     �D@      @      B@      ,@     �J@      =@      �?      @     �O@      T@      @      0@     �P@      @@     @T@     �J@     @Q@     @R@      @      (@     �N@     �Y@      &@      @     �a@      7@     �W@     �P@     @Y@     �W@      $@      (@     �I@      R@      &@      @     �[@      6@      J@     �H@      S@     @S@      $@              $@      >@              @      >@      �?      E@      1@      9@      2@              �?     �P@     �a@      (@      (@     �[@      ,@      u@      7@      t@     @T@      @              7@     �S@      @      @     �E@      @     �i@       @     @e@      A@                      &@     �C@      @      �?     �@@             �V@      @     @S@      2@                      (@      D@       @      @      $@      @      ]@      @     @W@      0@              �?     �E@     �O@      @      @      Q@      &@      `@      .@      c@     �G@      @      �?      @@     �L@       @      @     �M@      @     �[@      $@     �a@      D@      �?              &@      @      @              "@      @      2@      @      "@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJy�5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @{a`
�v@�	           ��@       	                    �?�5��7�@s           �@                           �?�V{�&x@�           �@                            �?�n^i@@�            0r@������������������������       ��Q]��c@3             T@������������������������       ������@�            `j@                          �;@R?u3�;@�            �u@������������������������       �3WQ[~U@�            0s@������������������������       �7&[�T@             F@
                           �?���Q�	@�           �@                          �4@k�P��	@�           d�@������������������������       �V��׳>	@�            �v@������������������������       ���
mt 
@�           h�@                            @�J��@           �z@������������������������       ��`a��@�            0r@������������������������       �����@R            �`@                          �4@e�b��O@B           �@                           @��B���@N           �@                           �?舩��� @�           P�@������������������������       ��7����?�            �p@������������������������       �"d$ �@            z@                           �?�BH�8@�            �n@������������������������       ����E@A            �Y@������������������������       ��D(m?B@\             b@                          �7@��L!E@�           (�@                           �?* =�lS@�            �w@������������������������       ��H��p�@|            �g@������������������������       ��%��z�@r            �g@                           �?�]�)}@           �z@������������������������       ����G@E            @\@������������������������       ���@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     0q@     ��@      ;@     �L@     P~@     �V@     ��@      m@     (�@     �t@      B@      9@     �h@      t@      2@      F@     �t@      Q@     w@     �g@     �v@      l@      ;@             �N@      X@       @      $@     @T@      @     �d@      ;@      a@      K@      @              ?@     �B@       @       @     �E@      @     @S@      2@      I@      2@      �?              @      @              @      *@      @      7@      @      3@                              <@      @@       @       @      >@      �?      K@      (@      ?@      2@      �?              >@     �M@               @      C@             �U@      "@     �U@      B@      @              6@     �G@              �?      @@              U@      @     �U@      <@      @               @      (@              �?      @              @      @      �?       @              9@     @a@     @l@      0@      A@      o@      O@     �i@     @d@     �l@     @e@      7@      9@     @[@     �b@      0@      :@     `h@     �H@     �`@     �Z@     `c@     @`@      5@      $@      6@      B@       @       @     @Q@      $@     �P@     �D@     �I@     �C@      "@      .@     �U@      \@      ,@      2@     �_@     �C@     �P@     @P@      Z@     �V@      (@              =@     �S@               @     �J@      *@      R@      L@     @R@      D@       @              3@      D@              @      H@      "@      F@     �B@      L@      >@       @              $@      C@               @      @      @      <@      3@      1@      $@              �?      S@     �n@      "@      *@     �c@      7@     0�@     �E@     �{@      Z@      "@             �D@     @^@      @      @     �G@      @     �y@      .@      n@     �D@       @              9@     @V@      �?      @      ;@      @     `t@      $@     �e@      7@                      *@      =@                      @             `b@       @      P@      @                      (@      N@      �?      @      6@      @     `f@       @     �[@      1@                      0@      @@       @       @      4@              U@      @     �P@      2@       @              @      0@              �?      @              D@      @      3@      @       @              "@      0@       @      �?      *@              F@             �G@      *@              �?     �A@     @_@      @       @     @[@      4@     �i@      <@     �h@     �O@      @              .@     �R@      @      �?      F@      (@     �Y@      @     @X@      2@      @              "@      E@      �?      �?      >@       @      E@             �G@      @      @              @     �@@      @              ,@      @      N@      @      I@      (@      @      �?      4@      I@      �?      @     @P@       @     �Y@      7@     �Y@     �F@      �?               @      2@                       @      @      F@      @      @@       @              �?      2@      @@      �?      @     �O@      @      M@      4@     �Q@     �B@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ7�chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�w�v@�	           ��@       	                    �?ޞ�D=�@
           x�@                           �?�}�hP@-           �}@                          �1@�]jg�"@s            �f@������������������������       ��W�_�0�?             B@������������������������       �(9x"&�@Z            `b@                          �<@&u0E@�            �r@������������������������       �K���@�            `o@������������������������       ��{Ԃ�V@            �F@
                            �?���dg@�           ��@                           @�p�(J(@{            �i@������������������������       �����k	@'            �Q@������������������������       �`���/s�?T            �`@                            @�4�G6�@b           ��@������������������������       � V>��@           �{@������������������������       �
v�h�" @N            �^@                          �8@��Ct�R@�           ֤@                          �1@��a�X@�           (�@                           @�a��@�            @w@������������������������       ��9K|^@k             f@������������������������       ���|)iq@�            �h@                            �?�rS�r�@�           X�@������������������������       �ܣľޝ@            {@������������������������       �`zd�@�           ��@                           �?��~���	@�           �@                          �;@2H{��
@�            `v@������������������������       ��j'lB	@o            �d@������������������������       �Ґ�g�:
@�             h@                          �<@3+	F��@�            �s@������������������������       �TP�}�,@�             k@������������������������       �7�BU�x@;            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      t@     �@      >@      H@     P{@     �V@     Ў@     @m@     ��@     �u@     �D@             �W@     �d@      @      $@      Y@      *@     �{@      G@     �q@     �T@      "@              H@     �R@      @      "@      G@       @     �Y@      @@     @Y@     �J@      @              2@      2@                      1@              K@      $@     �K@      $@      �?                      �?                      @              3@              $@                              2@      1@                      &@             �A@      $@     �F@      $@      �?              >@     �L@      @      "@      =@       @     �H@      6@      G@     �E@      @              ;@      J@      @      @      4@       @     �G@      1@      E@      <@      @              @      @               @      "@               @      @      @      .@                      G@     �V@              �?      K@      &@     u@      ,@     �f@      >@       @              @      ;@                      ,@      @      Z@       @     �C@      $@       @              @      @                      @      @      <@              3@      @       @                      4@                      $@      �?      S@       @      4@      @                     �E@     �O@              �?      D@      @      m@      (@     �a@      4@                      C@      M@                      =@      @     �e@      &@      [@      .@                      @      @              �?      &@             �M@      �?     �A@      @              2@     @l@     �w@      ;@      C@     u@     �S@     �@     �g@     ��@     �p@      @@      (@     `c@     0r@      &@      ;@     @n@      I@     �~@     �Z@     �z@     @d@      1@      �?      7@     �M@       @      @      3@       @      a@      4@      S@      >@              �?      3@      >@       @              &@       @      J@      0@      6@      5@                      @      =@              @       @              U@      @      K@      "@              &@     �`@      m@      "@      7@     �k@      H@     v@     �U@     0v@     �`@      1@             �H@     �H@      @      @      K@      "@      Z@      <@     �U@      C@       @      &@     �T@     �f@      @      2@      e@     �C@      o@     �M@     �p@     �W@      "@      @     �Q@     @U@      0@      &@     �W@      <@     �L@     @T@     @Z@     �Y@      .@      @     �B@      G@      .@      @     �F@      5@      7@      K@     �D@     �I@      .@              (@      4@       @              7@       @      (@     �A@      8@      (@      (@      @      9@      :@      @      @      6@      *@      &@      3@      1@     �C@      @              A@     �C@      �?      @      I@      @      A@      ;@      P@      J@                      2@      9@              @      8@      @      ?@      7@      K@     �@@                      0@      ,@      �?      @      :@       @      @      @      $@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�E{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�j�h�j@�	           ��@       	                    @�����@J           �@                          �1@{%a>m�@�           ��@                           �?c��9�@�            Pq@������������������������       �Ȑu�d@1             V@������������������������       �$]@�U@u            �g@                            @D=�gtU@            X�@������������������������       �Z��5�o@5           P�@������������������������       ��h'��@�            t@
                           �?��*ҹ�@�           ��@                           @��!���@l           ��@������������������������       �.F$~2@M             \@������������������������       ��ۚ��B@           @|@                          �1@��m���@8           �~@������������������������       ��X�O�6�?h            �d@������������������������       �U<7���@�            pt@                           �?"��>��@D           �@                            �?��?�	@-           �@                           @)�tI	@�            �o@������������������������       ��yU��S	@z            �f@������������������������       �9y�8�@/            @R@                          �?@m:
�Z	@�           �@������������������������       �����@d           x�@������������������������       ���ԏ�n@              J@                           @�e6F˿@           (�@                           �?z��ν�@�            �o@������������������������       �i�k�@(            �P@������������������������       �&w���E@r            �g@                           @�? >�@}           0�@������������������������       �)Ș2�@�            �y@������������������������       ��d�7 �@�             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     x�@      B@     �F@     P~@     �W@     ؏@      m@     �@     pv@      @@      @     �\@     @u@      .@      6@      n@      A@     ؅@     @V@     P{@     �d@      ,@      @     �T@     `h@      @      0@     �d@      4@     @n@     @R@     �h@      Z@      &@              5@      J@              @      ?@      �?     �T@      *@     �N@      *@                      @      $@                      (@      �?      B@       @      5@      @                      2@      E@              @      3@              G@      &@      D@      $@              @     �N@     �a@      @      *@     �`@      3@      d@      N@     @a@     �V@      &@       @     �E@      R@      @      @     �R@      &@      X@      F@     @Y@     �L@      "@      @      2@     �Q@      �?      @     �M@       @      P@      0@     �B@      A@       @             �@@      b@       @      @      S@      ,@     �|@      0@     �m@      O@      @              7@     �N@      @      @     �L@      &@     �m@      "@     �^@     �B@      �?              $@      4@                      @       @      B@      @      0@       @      �?              *@     �D@      @      @      I@      @      i@      @     �Z@      =@                      $@      U@      @      @      3@      @     �k@      @      ]@      9@       @                      0@                      @             @U@       @      I@      @      �?              $@      Q@      @      @      (@      @      a@      @     �P@      3@      �?      @     �f@     `k@      5@      7@     �n@     �N@      t@      b@     �r@      h@      2@      @     �X@     �^@      .@      0@     �b@      D@     �T@     @Y@     �\@     �Z@      ,@      �?      ?@     �@@      �?      "@     �E@      &@     �C@     �A@      <@      3@      @      �?      :@      9@               @      5@      "@      A@      1@      6@      .@      @              @       @      �?      �?      6@       @      @      2@      @      @      �?      @      Q@     �V@      ,@      @     @Z@      =@     �E@     �P@     �U@      V@      "@       @      K@     �U@      &@      @      X@      9@     �E@      P@     @T@      U@      "@      @      ,@      @      @      @      "@      @               @      @      @              �?     �T@      X@      @      @     @X@      5@     �m@     �E@     `g@     �U@      @              >@     �@@              �?      A@      &@     �K@      8@     �C@      :@       @              @       @                      @      �?     �@@       @      (@      @                      7@      ?@              �?      ;@      $@      6@      6@      ;@      7@       @      �?     �J@     �O@      @      @     �O@      $@     �f@      3@     �b@      N@       @      �?     �B@     �E@      �?              D@      @     `a@      "@      Z@      A@       @              0@      4@      @      @      7@      @      F@      $@      F@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJfwhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?9E���H@�	           ��@       	                   �5@�����@�           ��@                           �?:���N@m           ؁@                           �?jq�TK�@�            �j@������������������������       ���糩R@D            @Y@������������������������       �U�X�.@K            �\@                          �1@u�Z4 k@�            @v@������������������������       ����T0�?E            �[@������������������������       ���
�q@�            �n@
                          �8@	�Q4��@4           P~@                          �6@=��@�            �l@������������������������       ��OZ�q�@0            �Q@������������������������       ��o��5M@f             d@                           @6�Z+�I@�            �o@������������������������       �zzy��@e            �d@������������������������       ��V�@9             V@                           @���h@�           R�@                           �?֥ 4�@�           (�@                           �?��N��@           �|@������������������������       ��ٖX��@�             u@������������������������       ����{��@M             ^@                          �2@��~o�\	@�            �@������������������������       �3;)y�@�             j@������������������������       �%�+��	@           ��@                          �7@v�9��D@>           |�@                           @r#�@s�@w           ��@������������������������       ���&��@�           ��@������������������������       ��A�2�M@�            �p@                           @:�E��@�             t@������������������������       �8#%6C�@�            �p@������������������������       �����#�@            �K@�t�b��	     h�h5h8K ��h:��R�(KKKK��h��B�        *@     `s@     �@      8@      K@     P}@      U@     ��@     `l@     ؈@      w@     �A@       @     �Q@     `b@      @      0@     �\@      4@     0s@      R@     �i@      U@      $@              6@     �Q@              @     �H@      @      k@      @@     �_@     �C@      @              *@      9@              �?      >@      @     �D@      8@      K@      4@      @                      @              �?      4@       @      :@       @      ;@      $@                      *@      2@                      $@      �?      .@      0@      ;@      $@      @              "@      G@              @      3@      @      f@       @     @R@      3@                              (@              �?      @              R@       @      (@      "@                      "@      A@               @      0@      @      Z@      @     �N@      $@               @     �H@      S@      @      (@     �P@      ,@     �V@      D@      T@     �F@      @             �@@      7@      @       @     �A@      @     �M@      .@      ?@      .@       @              *@      "@      �?      @      @              ;@      @      @      @                      4@      ,@      @      @      ?@      @      @@      "@      <@      (@       @       @      0@     �J@              @      ?@      $@      ?@      9@     �H@      >@      @       @      (@      F@               @      6@      $@      0@      1@      ;@      .@                      @      "@               @      "@              .@       @      6@      .@      @      &@     �m@     �v@      3@      C@      v@      P@     H�@     `c@     `�@     �q@      9@      &@     �c@      j@      .@      <@     �m@      G@     �n@     @`@     �o@     @h@      4@             �L@      K@      @       @      P@      @     @[@      4@     �X@     �B@      @              G@      G@      @       @     �J@      @     �P@      0@      P@      =@      @              &@       @                      &@             �E@      @     �A@       @              &@      Y@     @c@      (@      4@     �e@     �E@      a@     �[@     �c@     �c@      0@       @      (@      5@       @      �?      8@             �K@      8@     �@@      @@       @      "@      V@     �`@      $@      3@     �b@     �E@     �T@     �U@     �^@     @_@      ,@             �T@     �c@      @      $@     �]@      2@     0}@      9@     �t@     �V@      @              I@     �^@       @      @     �Q@      (@      y@      *@     �o@     �L@       @             �A@     �S@      �?      �?      H@      @     �t@       @     `f@      A@      �?              .@     �F@      �?      @      6@      @     @R@      @     �R@      7@      �?              @@      B@       @      @      H@      @     @P@      (@     �S@     �@@      @              7@      <@              @     �A@      �?     �L@      &@     �R@      @@                      "@       @       @              *@      @       @      �?      @      �?      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{M�$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @A����T@�	           ��@       	                    �? %��-�@s           v�@                          �;@}oQ�f@�           P�@                          �1@��(x�l@`           ��@������������������������       �xC��& @A            @\@������������������������       ��P�+P�@           P|@                            �?�d�~@4             U@������������������������       ���1�@             1@������������������������       ����@)            �P@
                          �9@e��ho	@�           Ę@                          �3@�(��@�           h�@������������������������       ��S�(�k@            |@������������������������       �d�;�@�           І@                          �;@��e���	@�            py@������������������������       ��j`xq$	@^            @c@������������������������       �g�2��	@�            �o@                           �?5���@+           8�@                          �9@��W'o @g           ��@                           @�?Yes�?A           ��@������������������������       �N��)P�?�            v@������������������������       �=���� @n            �e@                           @X�ۂD@&             P@������������������������       �~ zdf�@            �@@������������������������       �/A�%� @             ?@                           @�h�ů>@�           ��@                          �2@����@           Ȉ@������������������������       ��W���
 @�             n@������������������������       �\��oD@`           H�@                          �4@ڵ��m@�            Pr@������������������������       ���r� �@N             ]@������������������������       ��fH{"=@q             f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@      r@     ��@      7@      K@     �|@     �S@     h�@     @l@     0�@     �u@     �@@      8@     �k@     Pu@      1@      F@     �t@     @P@     pw@      g@      w@     �m@      :@       @     �Q@     �V@      �?      $@     �T@      @      f@     �@@     �`@     �E@      @              N@     �S@      �?       @      Q@       @     �e@      6@     �^@      =@      @               @      3@                      2@              G@      @      4@      @                      M@     �M@      �?       @      I@       @     �_@      3@     �Y@      8@      @       @      $@      *@               @      ,@      �?      @      &@      (@      ,@       @       @      �?      @                      �?      �?                       @       @       @              "@      @               @      *@              @      &@      $@      (@              6@     �b@     @o@      0@      A@      o@      O@     �h@      c@     �m@     @h@      5@      $@     �Z@     `h@      (@      >@      i@      9@     �d@     �[@     �g@     �^@      ,@      @      ;@      N@      @      @     �P@      @      V@      K@     �R@      H@      @      @     �S@     �`@       @      7@     �`@      2@      S@      L@     �\@     �R@       @      (@     �F@     �K@      @      @      H@     �B@     �A@      E@      G@      R@      @              0@      2@       @              3@      0@      .@      9@      (@      9@      @      (@      =@     �B@       @      @      =@      5@      4@      1@      A@     �G@      �?       @     �P@     �o@      @      $@     ``@      *@     ��@     �D@     @y@      \@      @              *@     �W@               @      7@      @     Pr@      @     @a@      3@                      *@     �U@               @      4@      �?     @q@       @      ]@      &@                      "@      L@                      "@      �?     �h@             �R@      @                      @      ?@               @      &@             �S@       @      E@      @                               @                      @      @      1@      @      6@       @                              @                       @       @      &@              @      @                               @                      �?      �?      @      @      0@       @               @      K@      d@      @       @      [@      "@     u@      B@     �p@     @W@      @       @     �B@      \@      �?      @     �R@      @      q@      3@     `i@     �M@      @              @     �B@                      @             �Z@      @      Q@      0@               @      @@     �R@      �?      @     �Q@      @     �d@      0@     �`@     �E@      @              1@      H@      @      @      A@      @     �O@      1@     �O@      A@       @              @      5@      @       @      &@             �B@      �?      9@      &@                      (@      ;@       @      @      7@      @      :@      0@      C@      7@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ#<�vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�0DLm@�	           ��@       	                    @�����@�           ��@                           �?��`�@i           T�@                           �?T�uI=z@           Pz@������������������������       ��q[z�@�            0r@������������������������       ���	��@O            @`@                            �?Z��|w1	@]           ��@������������������������       �� *�Z	@+           �|@������������������������       ��o<V	@2           @~@
                            �?.$x�X@�           $�@                           �?��V�@           �x@������������������������       �QKC��$@�             k@������������������������       ��}&{&�@            �f@                           �?�/=GP�@�           ��@������������������������       �	��4>@�            �u@������������������������       �ߺVR��@�            �@                          �<@���ks]@�           ��@                           �?�1�e�@y           `�@                          �7@��'D@�            Pq@������������������������       �/*��Qp@�            �i@������������������������       �[�r$bg@-            �Q@                           �?w�k�)�@�           ��@������������������������       ���P�4	@           0{@������������������������       �𷥽��@�            @r@                          �=@�kt�@O            �_@                           �?Z���@             <@������������������������       ��D=�U�@             (@������������������������       �+�%W�@
             0@                          �>@'�E`�z@=            �X@������������������������       ���>�kk@             B@������������������������       �uO�[�@)            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     `r@     Ѐ@      6@      H@     �~@      X@     x�@     `j@     ��@     px@      B@      @      i@     px@      &@      B@     �t@     �N@     ��@     @b@      �@     pp@      7@      @     @`@      g@       @      <@      h@     �D@     �l@     �Y@      p@     �d@      5@      �?      G@      C@              @     �I@      @     @W@      2@      ]@      E@      @      �?     �@@      ?@              @     �C@       @     �K@      .@      Q@     �C@      @              *@      @              �?      (@      @      C@      @      H@      @       @      @      U@     `b@       @      8@     �a@      B@     �`@     @U@     �a@     �^@      ,@             �G@     @R@      @      ,@     @R@      *@     �R@      D@     �M@     �I@      &@      @     �B@     �R@      @      $@      Q@      7@      N@     �F@     �T@      R@      @             �Q@     �i@      @       @     @a@      4@     �@     �E@      t@     �X@       @              1@      C@      �?             �@@      @     `e@      *@     �U@     �@@                       @      2@                      .@      �?      X@      @     �I@      4@                      "@      4@      �?              2@      @     �R@      @      B@      *@                     �J@      e@       @       @     @Z@      0@      u@      >@     `m@     @P@       @              ,@     @P@                      3@       @     �`@      @     �U@      ,@       @             �C@     �Y@       @       @     �U@      ,@      i@      8@     �b@     �I@              .@     �W@     `b@      &@      (@      d@     �A@      n@     @P@     `j@      `@      *@      &@     @S@     �_@       @      $@     @`@      <@     @m@      L@     `i@     �Z@      *@              4@      8@                      .@      @     @[@      *@     �Q@      6@                      *@      *@                      @      @      V@      @     �O@      0@                      @      &@                       @              5@      $@       @      @              &@     �L@     �Y@       @      $@     �\@      9@     @_@     �E@     �`@     @U@      *@      &@     �B@      J@      @      @      W@      2@     �F@     �@@     �R@      K@      (@              4@     �I@      @      @      7@      @      T@      $@      M@      ?@      �?      @      1@      4@      @       @      >@      @      @      "@       @      5@                      @      @      �?              @      @              @      @       @                      @      �?                       @                      �?      @       @                      @       @      �?              �?      @              @                              @      &@      1@       @       @      ;@       @      @      @      @      3@                      @      @              �?      0@       @      @      �?              @              @       @      (@       @      �?      &@              @      @      @      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�%XGhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���[@�	           ��@       	                    �?�����@\           :�@                          �8@�mD%f�@�           ��@                           �?�Tg�@-           �~@������������������������       �@�p��@�            �h@������������������������       ���*^�@�            @r@                           �?�e�<�}@j            `e@������������������������       ��&�@@             �J@������������������������       �����@J            �]@
                           �?�'4$�	@�           (�@                           �?L����	@�           ̑@������������������������       �g�uO�D@6            �V@������������������������       ��� N�	@�           d�@                          �3@�X�zX@           py@������������������������       �:�1Y@^            @`@������������������������       �$�����@�            Pq@                            �?���l%@3           ��@                          �4@\/Vv�L@\           ��@                          �0@���[M@R           �@������������������������       �j��\���?%             O@������������������������       �+��%d@-           P~@                            �?��dt�@
           �y@������������������������       �jnN�x�@n            �c@������������������������       ��m�t�G@�            �o@                           @��2)�@�           h�@                          �3@5�����@M           ��@������������������������       ���x6!�?�            �l@������������������������       �'��@�            0s@                          �5@�aW��%@�            �j@������������������������       ���:��@@            �W@������������������������       ��W�-@J            �]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     X�@      ?@     �M@     @|@      U@     H�@      h@     p�@     �v@      C@      5@      j@     @v@      8@     �C@     t@      M@     pw@      d@      w@     `n@      >@             �M@     �^@      @      @      S@      @      d@      5@      b@     �O@      @              E@      T@      @      @      H@      @      a@      "@     �^@      D@      �?              1@      >@      @      @      5@      @     @Q@      @      >@      *@      �?              9@      I@                      ;@              Q@      @      W@      ;@                      1@      E@              �?      <@              7@      (@      7@      7@       @              @      &@                      &@              &@              @       @                      $@      ?@              �?      1@              (@      (@      2@      .@       @      5@     �b@     @m@      5@     �A@     �n@     �K@     �j@     �a@     �k@     �f@      ;@      5@     @]@      d@      1@      5@     `f@      E@     �b@     �Z@     `c@     �b@      9@      @      1@      @                      7@      @      @      "@      ,@      $@      �?      ,@      Y@     �c@      1@      5@     �c@     �C@      b@     @X@     �a@     @a@      8@             �@@     �R@      @      ,@     �P@      *@     �P@      A@      Q@      @@       @              @      @@               @      0@       @     �A@      (@      5@      @                      <@      E@      @      (@      I@      &@      @@      6@     �G@      ;@       @      �?     �U@     �l@      @      4@     ``@      :@     ؄@      ?@     �w@     @]@       @             �D@     ``@      @      (@     �T@      5@     �v@      2@     �j@     @Q@      @              1@      M@       @       @      D@      �?     �n@      @     �_@     �E@                              $@                                      >@              "@      *@                      1@      H@       @       @      D@      �?     �j@      @     �]@      >@                      8@     @R@      �?      @     �E@      4@     @^@      &@     �U@      :@      @              &@      3@      �?              *@      @      J@      @     �C@      ,@                      *@      K@              @      >@      ,@     @Q@       @     �G@      (@      @      �?      G@      Y@      @       @      H@      @     �r@      *@      e@      H@      @      �?      <@      M@               @     �B@      @     �n@      @     �`@      5@      �?              @      ?@              �?      @              a@      @      B@      @              �?      5@      ;@              �?      >@      @      [@       @     �X@      .@      �?              2@      E@      @      @      &@       @     �L@       @     �A@      ;@      @              (@      (@              �?      @      �?      C@       @      *@      "@      @              @      >@      @      @       @      �?      3@      @      6@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJj�:AhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�O��-@�	           ��@       	                    �?��=F�@U           
�@                            �?Y�)�	�@�           ��@                           �?�<X�@�            �i@������������������������       �|�_�	&@(            �N@������������������������       �����b&@\             b@                           �?l�1v��@S           X�@������������������������       ��iGo@�             m@������������������������       ��x_}y�@�            0r@
                           �??*����@~           ��@                          �3@�
z#p@N           8�@������������������������       ��er����?�            �x@������������������������       ��F���I@a             c@                           @���W��@0           0�@������������������������       ����j�@�            �y@������������������������       �q���@5           �~@                           @��(��@^           �@                           �?��71�M	@�           ��@                          �:@���HC�	@&           �@������������������������       ����4L	@Z           ��@������������������������       ����H�o	@�            Pt@                            �?O���@�            Pp@������������������������       ���L{F@-            @R@������������������������       ��nF�l�@u            �g@                           �?�qm��@�           ��@                            @CM��Q�@�            �s@������������������������       ���7o:@�            �o@������������������������       ���r�D� @$             N@                           @����@�            Pr@������������������������       ���a�4@�            �q@������������������������       �4S����?             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     h�@      7@     �L@      }@     �S@     �@     �m@     ȉ@     pt@      =@      @     �]@     r@       @      8@     @l@     �A@     �@      X@     �@     �c@      $@      @      N@     �V@      @      ,@     �\@      2@     @a@      H@     @d@     �P@      @              3@      ;@                     �B@       @     �@@      .@      N@      &@      �?               @      *@                      @              (@      �?      ;@      @                      1@      ,@                      A@       @      5@      ,@     �@@       @      �?      @     �D@     �O@      @      ,@     �S@      0@     @Z@     �@@     �Y@      L@      @       @      ,@     �B@      �?      @      6@      @     �K@      4@      H@      8@       @      @      ;@      :@       @      $@      L@      *@      I@      *@      K@      @@      @             �M@     �h@      @      $@     �[@      1@     ȁ@      H@     pu@     @V@      @              8@      P@              @      @@      @     Pq@      $@     �]@      4@                      5@      @@                      .@             �i@      @      Y@      0@                      @      @@              @      1@      @     �Q@      @      2@      @                     �A@     �`@      @      @     �S@      ,@     @r@      C@      l@     @Q@      @              0@     �T@       @             �G@      "@     @]@      =@     �Q@     �A@      �?              3@      J@      @      @      @@      @     �e@      "@     `c@      A@       @      (@      g@     �m@      .@     �@@     �m@     �E@     �s@     �a@      t@     `e@      3@      &@      a@     �b@      "@      9@     �e@      B@     @b@     �]@      e@     �`@      0@      &@     @\@      ]@      "@      2@     ``@      >@     @W@     @W@     @_@      \@      ,@      @      T@     �T@      @      &@     �Q@      "@      O@      P@     �V@     �I@      (@      @     �@@      A@      @      @     �N@      5@      ?@      =@     �A@     �N@       @              8@     �A@              @     �E@      @     �J@      9@      F@      6@       @              @      &@              �?      (@       @      2@      @      &@      "@       @              4@      8@              @      ?@      @     �A@      6@     �@@      *@              �?     �G@     @U@      @       @      P@      @     �e@      8@     �b@     �B@      @      �?      >@      H@      �?      @      ?@      @     @W@      @     @R@      3@      @      �?      >@      C@      �?      @      ;@      @     @P@       @      N@      1@      @                      $@               @      @              <@      �?      *@       @                      1@     �B@      @       @     �@@       @      T@      5@     �S@      2@                      &@     �A@      @       @     �@@       @      T@      3@     �S@      2@                      @       @      �?                                       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��~�-@�	           ��@       	                   �1@���LB�@u           >�@                           �?lt�>@�            �q@                            �?�aAU��@6            �T@������������������������       �E�B{�@             C@������������������������       �\�6�\ @            �F@                           �?QW�%�@            �h@������������������������       ��13�7@=            �W@������������������������       ��%vl:@B            �Y@
                           �?�{`�	@�           �@                           �?/ގ�8)@C           @�@������������������������       ����t0�@�            �w@������������������������       ��ӿ�@Z             a@                          �9@5���s�	@}           ��@������������������������       �LW]lA	@           ��@������������������������       ����r޴	@�            �x@                          �5@�pr��@F           ��@                           �?'�|�G@�           �@                          �4@d�]��L�?�            y@������������������������       �l<�!���?�             u@������������������������       �^��)�?%            @P@                           �?'��>�w@�           P�@������������������������       �@,ɠB�@�            �t@������������������������       � qߌx�@�            �u@                           @��	Z�@�           x�@                           �?9Y�u�@           �z@������������������������       �f(��@�            �k@������������������������       �h���TL@�            �i@                           @��0��@}            `h@������������������������       �{ğ-5@r             f@������������������������       ����N�@             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     Ps@     �@      7@      J@      |@     @T@     X�@     �h@     ��@      v@      =@      5@     �i@     �t@      4@     �D@     @t@      O@      w@     �d@     �y@      m@      ;@      �?      "@     �K@                      :@       @      U@      (@      Q@      8@                      @      @                      @       @      =@      @      9@      @                       @      @                       @       @       @              (@      @                       @      �?                      @              5@      @      *@      �?              �?      @      H@                      4@             �K@      "@     �E@      1@              �?      @      >@                      .@              ,@       @      4@      "@                      �?      2@                      @             �D@      @      7@       @              4@     �h@     @q@      4@     �D@     �r@      N@     �q@     @c@     Pu@      j@      ;@      �?     �K@     �Q@      @      $@     �Q@       @     �\@      <@     �]@     �C@      @      �?      D@     �M@      @       @      K@      �?     �Q@      8@     �T@      A@      @              .@      (@               @      0@      �?      F@      @      B@      @       @      3@     �a@     �i@      .@      ?@     �l@      M@     @e@     �_@     �k@     @e@      5@      $@     �W@      c@      (@      7@     @f@      <@     @a@      T@      f@     �Y@      2@      "@     �G@      J@      @       @      I@      >@      @@      G@      G@      Q@      @              Z@     �n@      @      &@      _@      3@     ؂@      ?@     �{@     �]@       @             �J@      d@      �?      @      J@       @     �{@      ,@     0r@      J@       @              0@      O@              �?      @      �?     �k@      @     �S@      "@                      0@      D@              �?      @              h@      @     �P@      "@                              6@                      �?      �?      =@      �?      &@                             �B@     �X@      �?      @     �F@      @     �k@       @     �j@     �E@       @              4@      C@      �?       @      A@      @      [@      @      Z@      1@       @              1@      N@              @      &@      @     �\@      @     @[@      :@                     �I@     �U@       @      @      R@      &@      d@      1@      c@     �P@                      8@     �N@      �?      @     �D@      &@      `@      *@     @]@      <@                      1@      D@              @      9@       @     �Q@      @      G@      ,@                      @      5@      �?              0@      "@      M@      $@     �Q@      ,@                      ;@      9@      �?      �?      ?@              ?@      @      B@     �C@                      6@      8@              �?      9@              >@       @      A@     �C@                      @      �?      �?              @              �?       @       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJFWenhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@(�䁪@�	           ��@       	                    �?ZC����@:           x�@                          �1@��+ݦ@           x�@                          �0@^���+ @�             o@������������������������       ��o�.�4 @3            @T@������������������������       �$$z��p�?h            �d@                           @��1$u@�           ��@������������������������       �K��|B�@�            pr@������������������������       ���c<��?�             q@
                           @T|�|�@           4�@                           �?�>ޙ�@5           `�@������������������������       ��b?y��@�           x�@������������������������       ���$I�@�            �o@                          �5@G�_8:@�           �@������������������������       ����@�           h�@������������������������       �B.�F�@5             U@                          �<@��sǛ�@w           4�@                           �?���QF@�           8�@                          �9@��}��l	@F           p�@������������������������       �^�)R�@�            �s@������������������������       ��*�$�	@�            `j@                           @$iiEG@d            �@������������������������       �����Ks@/           P~@������������������������       �Z
3��@5            �V@                           �?�y����@�            �s@                           �?O
��*�@7            �U@������������������������       ��:�}.�@             E@������������������������       �	(0,�@            �F@                            @Y)�	@�             m@������������������������       ��iWx�B@]            �b@������������������������       ��x�v#	@9             U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@      r@     ��@      :@     �J@     �|@     �T@     H�@     �k@     ��@      v@      7@      $@     `c@     �v@      *@      :@     �o@      ?@     x�@     @_@     `�@     �d@      @             �F@     �[@              �?      M@      @     �u@      7@     @g@      B@      �?              *@      9@                      .@             �`@      @     �F@      &@                       @       @                       @              E@              ,@      @                      &@      1@                      @             @W@      @      ?@      @                      @@     �U@              �?     �E@      @     �j@      3@     �a@      9@      �?              ?@      F@              �?      A@      @     �S@      ,@      Q@      3@      �?              �?      E@                      "@      @     �`@      @     @R@      @              $@     �[@      p@      *@      9@     @h@      8@     @{@     �Y@      w@     ``@      @      $@     �T@     �b@      @      2@     �a@      2@      c@      V@     �b@     �U@      @      $@     �P@     �[@      @      .@     �X@      ,@     �T@     �P@      ]@     �P@      @              .@      C@      @      @     �F@      @     @Q@      6@      A@      4@                      <@      [@      @      @     �I@      @     �q@      ,@     �k@      F@      �?              6@     �W@      @      @     �D@      @     �n@      ,@     `j@     �C@      �?              @      *@      @              $@              C@              "@      @              @     �`@     �e@      *@      ;@     �i@      J@     @k@     @X@     Pr@     `g@      0@      @      Y@     �`@       @      5@     �c@     �A@     �f@      T@     @o@     �]@      (@       @      M@     @Q@       @      .@     @X@      7@     �I@      G@     @V@      M@      $@              D@     �F@      @      (@      R@      $@      4@      1@      K@     �@@      @       @      2@      8@      @      @      9@      *@      ?@      =@     �A@      9@      @      �?      E@     �P@              @     �M@      (@     �`@      A@      d@     �N@       @      �?      6@      J@              @     �J@      $@     @^@      3@     `b@     �J@      �?              4@      ,@                      @       @      &@      .@      ,@       @      �?             �@@      D@      @      @     �I@      1@     �A@      1@     �E@      Q@      @              @      ,@              �?      $@              0@      @      .@      6@      �?              �?       @              �?      �?              @      @      @      .@                      @      @                      "@              $@      �?       @      @      �?              =@      :@      @      @     �D@      1@      3@      *@      <@      G@      @              ,@      "@      �?      �?     �A@      "@      "@      "@      5@     �B@      @              .@      1@      @      @      @       @      $@      @      @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @V@��_@�	           ��@       	                    @�B���@           ��@                           �?e6�u��@h           P�@                          �<@��זLV@�            �x@������������������������       �@.3�@�            �u@������������������������       �d��t�@             G@                           �?��4�G	@i           H�@������������������������       �F�5
�L	@&            �L@������������������������       �A���	@C           ��@
                          �6@5(���@�           ��@                           @5��'dP@�           h�@������������������������       ������@`           ��@������������������������       ���ڀ�,@@           �~@                           �?p�<��@�             y@������������������������       �L9Xd�^@             j@������������������������       �1_�K�<@~             h@                           �?�Y{��2@�           ,�@                          �<@ť���@�            @s@                           �?B�T�@�            �q@������������������������       �b� j@_            �b@������������������������       ��W�j�o�?U            �`@������������������������       �֮!�0@             9@                           �?�#�$��@�           ��@                           @9��)X	@�            ps@������������������������       ��,e�2	@�            �q@������������������������       �z>�@             8@                           �?��.|�@3            ~@������������������������       �H_PhG�@!            �I@������������������������       �dƞ�*@           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        7@      r@     ��@      >@     �Q@     �|@     @T@     8�@      m@     ��@     @u@      8@      @      j@     0z@      3@     �F@     Ps@     �I@     h�@     �e@     8�@     @m@      1@      @      a@      j@      ,@      >@     �g@     �C@     @m@     �a@     �k@     �`@      "@             �H@     �H@      �?      @     �E@      @      Y@      8@     �U@      A@      �?             �B@      D@      �?      @      C@      @      Y@      5@     @T@      7@      �?              (@      "@                      @                      @      @      &@              @      V@      d@      *@      ;@      b@     �A@     �`@     @]@     �`@     @Y@       @      �?      @      @              @      $@      @      �?      &@      @      @       @      @     �T@     �c@      *@      5@     �`@      ?@     �`@     �Z@     �_@     �W@      @              R@     @j@      @      .@     @^@      (@     �@      ?@     �t@     �X@       @             �@@     @c@      @      &@     �P@      "@     }@       @     �m@     �M@      @              5@     �T@       @              @@      @     �q@      @     @Y@      >@                      (@      R@       @      &@      A@      @     �f@      @      a@      =@      @             �C@      L@      �?      @     �K@      @     �T@      7@      W@      D@      @              :@      E@              @      <@             �D@      @     �D@      1@      @              *@      ,@      �?      �?      ;@      @     �D@      2@     �I@      7@              0@     @T@     �a@      &@      :@     �b@      >@     p@      N@     �j@     �Z@      @              9@      ;@      �?      @      @@       @     �Y@      ,@      T@      2@                      9@      :@      �?       @      :@       @      Y@      &@      S@      ,@                      3@      6@      �?       @      &@       @      E@      $@      <@      (@                      @      @                      .@              M@      �?      H@       @                              �?              @      @               @      @      @      @              0@      L@     �\@      $@      3@      ]@      <@     `c@      G@     �`@      V@      @      "@      .@      F@      @      @     �D@      3@     �K@      &@      L@      G@       @      @      .@      C@      @      @     �@@      3@      K@      &@     �K@     �D@       @      @              @                       @              �?              �?      @              @     �D@     �Q@      @      *@     �R@      "@      Y@     �A@     �S@      E@      @       @      @      @              @      .@       @      @      @      @      �?              @      A@     �P@      @      "@      N@      @     �W@      <@      S@     �D@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ)e�_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����o�@�	           ��@       	                    �?���	@            T�@                            �?S{`Ur@+           �}@                           �?��emF@W            �]@������������������������       �������@$             J@������������������������       �l���@3            �P@                            @�����7@�            `v@������������������������       �끁�)@X            �d@������������������������       ����n��@|            @h@
                           �?�C�M�	@�           ��@                           @�SZ�_r@           �z@������������������������       �U��q��@I            �]@������������������������       �p�	H��@�            `s@                          �8@[!{�B
@�           `�@������������������������       �X��g�n	@           pz@������������������������       ��[Ո�g
@�            Pr@                          �4@:G�6��@�           �@                            �?��'s@�           T�@                           �?��~@�            0r@������������������������       ��!˫d�@U            �`@������������������������       ���r}P�?^            �c@                           @
m0K��@:           ��@������������������������       �z�#�A@           `z@������������������������       ��Mܴ�H@+           �|@                           @H��nN@�           |�@                           @D�9@�           �@������������������������       �)�g��@�            �s@������������������������       �X��|�^@�             x@                          �?@�1�	�@            z@������������������������       ��[C��_@           �x@������������������������       �ð]b�P@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �t@     ��@      B@     �G@     �|@     @T@     ��@     �m@     ��@     �s@      C@      6@     `h@     �k@      >@      ;@     p@     �E@     �i@     �b@     �o@     @g@      =@       @      L@     �P@      @      @      P@      �?     @V@      >@     @Z@     �G@      @       @      (@      9@                      @      �?      5@      @      A@      @      @       @      @      *@                      @      �?       @      @      .@       @                       @      (@                      @              *@      @      3@      @      @              F@      E@      @      @     �L@              Q@      8@     �Q@      D@       @              2@      4@      @       @      ?@              4@       @      C@      6@       @              :@      6@      @       @      :@              H@      0@     �@@      2@              4@     `a@     @c@      8@      7@      h@      E@     �]@     @^@     �b@     `a@      7@      @     �A@      P@       @      (@      T@       @     �Q@      =@     �N@     �M@      @      @      @      ,@       @      �?      8@      @      ,@      1@      2@      .@       @              >@      I@              &@      L@      @      L@      (@     �E@      F@      @      1@      Z@     �V@      6@      &@     @\@      A@      H@      W@     �U@      T@      2@      @      O@     �M@      @       @     @S@      .@      :@      A@     @Q@     �H@      $@      $@      E@      ?@      .@      @      B@      3@      6@      M@      2@      ?@       @             `a@     �u@      @      4@      i@      C@     �@      V@     �@     @`@      "@              P@     �e@      @      "@     @P@      @     �}@      @@     �q@     �M@      �?              $@     �@@               @      4@      �?     �b@      @     �K@      ,@                      @      (@               @      2@              K@      @      @@      "@                      @      5@                       @      �?      X@      @      7@      @                      K@     �a@      @      @     �F@      @     �t@      :@      l@     �F@      �?              A@      H@              @      1@       @      f@      2@     �X@      5@      �?              4@     @W@      @      �?      <@      @      c@       @     �_@      8@                     �R@     `e@       @      &@      a@      ?@     @r@      L@     �p@     �Q@       @             �K@      U@               @     �U@      8@     �i@      A@      d@      C@      @              @@      I@              @      C@      ,@     @P@      9@     �O@      4@       @              7@      A@               @      H@      $@     �a@      "@     @X@      2@      @              4@     �U@       @      @      I@      @     �U@      6@     �Z@     �@@      �?              1@     �U@       @      @     �G@      @     �U@      1@     �Y@      <@      �?              @                              @      @              @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�\8F@�	           ��@       	                    @��H致@           �@                            �?�V"P�@�           Ȅ@                          �;@�����b@�            �i@������������������������       �݇�0ߛ@w            �g@������������������������       �XL��J@
             *@                            �?Hb	ٕ�@&           �|@������������������������       �lbI8��@o            `e@������������������������       �U�@�             r@
                           @"��A]@a           �@                          �4@;��.���?�            �u@������������������������       �����T��?�             n@������������������������       �_�z> �@M            �[@                           �?�:<g�@u            `h@������������������������       �9r;'�8@;            �X@������������������������       �D�"=	r@:            @X@                           �?AJ�k4@�           �@                          �5@�Z��c�@�            �j@                          �1@� j@F            �[@������������������������       ��i�7��@
             3@������������������������       ��BeM1@<             W@                          �7@ű\�@A            @Y@������������������������       ���@             ;@������������������������       �d��7�@-            �R@                            �?k�.N�@H           v�@                           @Z���@�           �@������������������������       �S`nTYm@w           ��@������������������������       �`��F� 	@A            @Y@                          �1@�r�Dީ@�           ��@������������������������       �S;��z@�            q@������������������������       ���k�@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �t@      �@      6@     �H@     �}@     @V@     ��@     `i@      �@     �v@      >@             �V@     `d@       @      (@     �[@      (@     z@      =@     �q@     @U@      @             @R@     �U@       @      $@     �S@       @     �d@      9@     �b@      M@      @              2@      ?@              @      *@      @      H@      @     @P@      ,@       @              0@      ;@              @      (@       @      H@      @     @P@      &@      �?               @      @                      �?       @                              @      �?             �K@      L@       @      @     �P@      @     �]@      3@     �U@      F@      @              5@      2@       @      �?      5@              E@      $@      ?@      6@      @              A@      C@              @     �F@      @     @S@      "@     �K@      6@                      2@      S@               @      ?@      @     @o@      @     �`@      ;@      �?              ,@     �F@                      0@      @      g@             �S@      "@                      &@      6@                      $@              a@             �L@      @                      @      7@                      @      @      H@              5@      @                      @      ?@               @      .@      �?     @P@      @      K@      2@      �?              @      2@               @       @      �?      C@              1@      &@                      �?      *@                      @              ;@      @     �B@      @      �?      .@     `n@     �w@      4@     �B@      w@     @S@     ��@     �e@     H�@     �q@      8@      @      5@      ;@               @     �F@      .@      ,@      8@      =@      9@                      @      0@              @      7@      @      &@      $@      5@      1@                                                      @              @      @       @      @                      @      0@              @      4@      @      @      @      3@      (@              @      1@      &@              @      6@      "@      @      ,@       @       @               @      @      @              �?      �?      @      @       @      @      �?               @      &@       @              @      5@      @              (@      @      @              &@     �k@      v@      4@      =@     0t@      O@     (�@     �b@     �~@     �o@      8@             �P@      U@      @      @     �X@      3@     �d@      M@     �]@     �O@      ,@             �L@     �Q@      @      @     �W@      (@     �b@      G@     �Z@      F@      "@              $@      *@      �?      �?      @      @      1@      (@      (@      3@      @      &@     `c@     �p@      .@      6@      l@     �E@     �w@      W@     Pw@      h@      $@      �?      ,@     �A@               @      1@             @W@      @     �S@      :@              $@     �a@     `m@      .@      4@      j@     �E@     r@     @U@     pr@     �d@      $@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJqD5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�,��@�	           ��@       	                    �?8p]��n@M           Ġ@                            �?�[`9k@�           ȇ@                           @�0�@            �i@������������������������       ���_��@E            �[@������������������������       ��>�V��?:             X@                           �?�+ҵ�@R           P�@������������������������       �5L�BY@�            �q@������������������������       �V� Õ@�            �p@
                           @�����@|           ��@                          �2@A��@�           ��@������������������������       �s��l_@�            �r@������������������������       �<��4"	@           0z@                           @M��9�@�           Ȅ@������������������������       ���]
�@�            �q@������������������������       ��-��l@�            �w@                            �?e<:��@f           ��@                          �<@o���@e           ��@                           @��Mm�@�           ��@������������������������       ��(4���@�           (�@������������������������       ��Y9D�@             :@                           @§�֮>@s            �f@������������������������       �03֛�@P            �]@������������������������       �2�Bf�@#            �O@                           �?y��J�@           ��@                           �?��m@�            �k@������������������������       �㆓	k@=            @W@������������������������       �W�KH!�@P             `@                          @@@����>@t           ��@������������������������       �/d��*@f           ��@������������������������       �.�h�M@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     ��@      @@     �I@     �z@      S@     ��@     �i@     �@     @v@      ?@      @     @\@     @s@      0@      5@     �h@      7@     (�@     @W@     �~@     �d@      $@              F@     @W@               @     �F@             �s@      3@      h@      F@      @              @      >@              �?      *@              V@      �?      L@      ,@                      @      7@              �?       @              ;@      �?      D@      @                              @                      @             �N@              0@      @                      D@     �O@              �?      @@             �l@      2@      a@      >@      @              0@      ?@                      ,@             �`@      ,@     �L@      1@      @              8@      @@              �?      2@              X@      @      T@      *@              @     @Q@     �j@      0@      3@     �b@      7@     px@     �R@     pr@      ^@      @      @      H@     �_@      *@      (@      [@      0@     �^@      Q@     @^@     �R@      @      �?      4@     �F@              @     �I@      @      Q@      @@     �E@     �@@      �?      @      <@     @T@      *@      "@     �L@      (@      K@      B@     �S@      E@      @              5@     @V@      @      @     �E@      @     �p@      @     �e@     �F@      �?               @     �I@       @              6@      @     @X@      @     �P@      9@                      *@      C@      �?      @      5@      �?     �e@      �?     �Z@      4@      �?      $@     `g@     �o@      0@      >@     `m@     �J@     �s@     �[@     �u@      h@      5@       @     @[@      _@      &@      2@     �]@     �B@     �c@      R@     �h@     @]@      *@       @     �U@     @W@      &@      .@     �Z@      :@     @b@      O@     `e@     @P@      "@       @      U@     �V@      $@      .@     �Y@      7@     @b@     �I@     @e@      P@       @               @       @      �?              @      @              &@      �?      �?      �?              7@      ?@              @      &@      &@      $@      $@      :@      J@      @              *@      0@              @      @      $@      @       @      *@      E@      @              $@      .@                      @      �?      @       @      *@      $@               @     �S@      `@      @      (@     @]@      0@     �c@     �C@     �b@     �R@       @              5@      D@      �?      @      5@       @     �P@       @      G@      *@                      $@      :@      �?      @      .@              (@      @      .@      @                      &@      ,@                      @       @      K@      @      ?@      @               @     �L@      V@      @      "@      X@      ,@      W@      ?@     �Y@      O@       @      �?     �H@      V@      @      "@     �W@      ,@      W@      =@      Y@      J@       @      �?       @                               @                       @      @      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJձ�ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @�QR�f.@�	           ��@                          �3@�o�Y�@}           R�@                           @/d䭬v@�           x�@                           @ʁ<�@�            �@������������������������       �8ʧ�#�@h           ȁ@������������������������       ��7����@U            `a@������������������������       �)��B�N@             &@                          �;@�15�H	@�           h�@	       
                   �7@H�����@�           ��@������������������������       �i��cp@�           ��@������������������������       �Ĕ�}�@(           @}@                           @5o��E�	@�             s@������������������������       ��-j�r|
@�             j@������������������������       �t�[�@5             X@                          �1@n��h_�@:           ��@                           �?}+-.͠�?�            �v@                           @�Q�{���?{            �g@������������������������       ����5�?d            �c@������������������������       ��(Ռ��?             >@                           @!Ԋ����?f            �e@������������������������       �������?0             S@������������������������       ����:��?6            �X@                           �?~QF;
�@Y           Д@                            @lL̐�@           �y@������������������������       ��0- �"@�            �u@������������������������       ���� �?,             Q@                           @���3C�@X           ��@������������������������       �m�F��@�           @�@������������������������       �^􁔪@Y            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@      q@      �@      :@      K@     P|@     �U@     T�@     �j@     h�@      v@      =@      4@     �f@     �u@      3@      D@     @t@     �P@     �x@     �f@     @w@      n@      7@      @      K@     @\@      @      �?      S@       @     �i@      M@     @`@      N@      @      @      K@      \@      @      �?     �R@      @     �i@      M@      `@      N@              @      D@     �U@      �?      �?      M@      @     �d@     �A@     �]@      J@                      ,@      9@      @              1@             �C@      7@      $@       @              �?              �?                      �?       @      �?               @              @      .@      `@     @m@      .@     �C@      o@     �M@      h@     @_@     @n@     �f@      4@      @     �X@     �h@      $@      <@      k@      E@     �d@     �V@     �i@     �\@      1@      @     �Q@     @^@      @      2@     @a@      4@     �Z@     �E@      `@     �N@      "@              <@      S@      @      $@     �S@      6@     �M@      H@     @S@      K@       @       @      >@     �B@      @      &@      ?@      1@      ;@      A@      B@     @P@      @      @      9@      =@      @       @      5@      *@      0@      1@      9@     �C@      @      �?      @       @              @      $@      @      &@      1@      &@      :@                     �V@     �l@      @      ,@      `@      3@     0�@      @@     �y@     �\@      @               @     �F@              @      .@             �g@       @     �U@      (@      �?               @      <@              @      @             @Z@              B@       @                       @      8@              �?      @              V@              @@       @                              @              @      �?              1@              @                                      1@                      $@             @U@       @      I@      $@      �?                      @                      @              H@      �?      &@      @      �?                      (@                      @             �B@      �?     �C@      @                     �T@      g@      @      "@     �\@      3@     �|@      >@     0t@     �Y@      @              .@     �M@      �?       @      2@      @     �g@      @     �Y@      ,@                      (@      L@      �?              1@      @     �a@      @     @V@      ,@                      @      @               @      �?             �F@              ,@                              Q@     @_@      @      @      X@      *@     �p@      7@     �k@      V@      @             �F@     @[@      @      @      U@      "@     �m@      .@     �g@     �R@      �?              7@      0@       @              (@      @      =@       @      ?@      ,@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ,PrhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @���G9l@�	           ��@       	                     �?��G�@l           V�@                           �?�i���@�           ��@                           �?�h�Ol@|            �i@������������������������       �Uʈ[�j@0            �Q@������������������������       ����Ȧ@L             a@                          �1@dˣ��j	@!           �|@������������������������       ����fN@            �K@������������������������       �=�q�	@           py@
                          �<@�C�M��@�           <�@                          �5@��G�`@h           p�@������������������������       ��S�@�           P�@������������������������       �]X�ֹ�@�           ��@                            �?(K��@g            `f@������������������������       �����]@            �I@������������������������       �-@I@�@L             `@                           @���]m\@,           x�@                           �?`;k��@�           ��@                          �9@��*�@V           h�@������������������������       ��X<�@5           �~@������������������������       ��s���@!            �P@                           �?���.�@t           ��@������������������������       �6���^�@)            �M@������������������������       ��?�H@K           ��@                          �;@�#qv@b             d@                          �3@�ۗ{b�@V            �a@������������������������       ��'E��@#             O@������������������������       �'2�m0q@3             T@������������������������       ����r�?             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        :@     Ps@      �@      <@     �L@      ~@      S@     ��@     @h@     H�@     �v@     �E@      9@     @k@     Pt@      3@     �C@     �u@      L@     Pw@     `c@     0x@     �m@     �A@      @     �Q@     @V@      @      "@     �^@      5@     �]@     �I@     �Z@      K@      2@      @      1@      <@               @     �H@       @     �H@      &@      =@      0@              @      @      &@                      <@       @      (@      @      @      �?                      (@      1@               @      5@             �B@      @      :@      .@              @     �J@     �N@      @      @     @R@      3@     @Q@      D@     @S@      C@      2@              @      ,@                       @              "@      &@      .@      �?              @      I@     �G@      @      @     �Q@      3@      N@      =@      O@     �B@      2@      2@     �b@     �m@      0@      >@     `l@     �A@     �o@      Z@     �q@      g@      1@      (@     �^@     �i@      .@      :@     @i@      8@     @n@      U@      q@     `b@      1@      @      I@      ]@      @      3@     �[@      *@      d@      F@      e@     �S@      @       @     @R@     �V@      "@      @     �V@      &@     @T@      D@     @Z@     @Q@      $@      @      9@      >@      �?      @      9@      &@      *@      4@      @     �B@               @       @      @                              @      @      @       @      5@              @      1@      :@      �?      @      9@      @      "@      .@      @      0@              �?     �V@     �k@      "@      2@     �`@      4@      �@     �C@     `x@     �^@       @      �?      R@     �i@      @      2@     �\@      0@     ��@     �@@     �v@      [@       @              6@     �R@      �?      @      @@      @     �p@      $@      ]@      8@       @              6@      P@      �?      @      9@             �m@      $@      Z@      6@       @                      &@                      @      @      ;@              (@       @              �?      I@     @`@      @      .@     �T@      "@     �t@      7@     @o@      U@              �?      @      *@              �?      @      @       @      @      4@       @                      G@     @]@      @      ,@     �S@      @      t@      4@     �l@     �T@                      3@      2@      @              2@      @     �G@      @      8@      ,@      @              1@      2@      @              @      @     �G@      @      6@      &@      @              @      @                      @              <@              &@       @                      (@      (@      @              @      @      3@      @      &@      @      @               @                              &@                               @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�p!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @��}@�	           ��@       	                    �?���
�@�           ��@                           �?L2j,�6@�           �@                           �?�EC{�@�            �r@������������������������       �X�+K	@�            �k@������������������������       ��S��@4             S@                           �?E��l�@�            �u@������������������������       ��8���@�             o@������������������������       ��ҕ�@:            �W@
                           �?��
�A�	@�           �@                           �?�
�	@�           ��@������������������������       ��x��	@�            �v@������������������������       ���n�k	@�           ��@                          �4@/͒��@           �y@������������������������       �;���W@x            �h@������������������������       ��asݾ�@�            �j@                           @��;��!@           �@                           @�Z�d�%@�           �@                          �2@[�/|w@�             y@������������������������       ��F↘�?L            �^@������������������������       �����@�            �q@                           �?��Ę�&@�           ��@������������������������       �҇:�Д�?            �j@������������������������       �����Y@T           ؀@                          �>@�!��h�@R           �@                           �?�R��@@E           �~@������������������������       �ݵ�l�@            @g@������������������������       �r$��Em@�            �r@������������������������       ��#�Z�n@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     0r@     (�@      =@     @P@     �}@     �T@     ��@     �m@     �@     �x@      ;@      .@     �j@     t@      5@      J@     0u@      Q@     Pw@      h@     �v@     �p@      9@             �L@     @V@      �?      �?     @U@      @     �d@     �B@     �`@     �O@      @              9@      E@      �?      �?     �F@      @     @T@      4@     �J@      7@      �?              4@     �A@      �?      �?     �@@      @      I@      1@     �E@      0@      �?              @      @                      (@      �?      ?@      @      $@      @                      @@     �G@                      D@              U@      1@     @T@      D@      @              ;@      D@                     �@@             �D@      .@     �K@     �B@      �?              @      @                      @             �E@       @      :@      @       @      .@     `c@      m@      4@     �I@     �o@     �N@      j@     �c@     `l@     �i@      5@      .@     @_@     �c@      0@      @@     `i@     �F@     �`@     @\@     �d@     @d@      5@      "@     �E@     �J@      @       @     �S@      4@      9@      ?@      8@     �L@      @      @     �T@     @Z@      "@      8@     @_@      9@     @[@     �T@     �a@     @Z@      0@              >@     �R@      @      3@     �I@      0@     �R@     �E@      N@      E@                      @     �G@      @       @      4@      �?     �K@      .@      6@      6@                      9@      ;@              &@      ?@      .@      3@      <@      C@      4@              �?     �S@     �l@       @      *@     �`@      .@     �@     �F@     �y@      `@       @      �?     �L@     �b@              @     �T@       @     �|@      >@     �q@     @S@      �?      �?      @@     �M@               @      >@       @     �b@      *@     �T@      9@                       @      5@                       @             �Q@      @      &@      @              �?      8@      C@               @      <@       @     �S@       @      R@      4@                      9@     �V@              @     �J@             �s@      1@      i@      J@      �?              @      3@                      $@             @a@      �?      B@      @                      5@      R@              @     �E@             �e@      0@     �d@     �F@      �?              6@     �S@       @       @      I@      @      b@      .@     �_@     �I@      �?              0@      S@      @       @     �H@      @      b@      ,@     @_@      F@      �?              @      ;@      �?       @      "@             �T@      @     �E@      (@                      $@     �H@      @      @      D@      @     �N@      &@     �T@      @@      �?              @       @      @              �?      �?              �?      �?      @        �t�bub�{     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�E�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �5@*x�|_]@�	           ��@       	                    @�H�$�@_           "�@                           �?+��,�@�           X�@                           �?Q�7��@�            `w@������������������������       ���\��@r            `g@������������������������       ��6m-�@y            `g@                           �?'ݷ���@�            �@������������������������       ���>u-,	@F           �~@������������������������       ��=�O�F@�             n@
                           �?q5���@�           �@                           @=�l� @�             y@������������������������       �^�c�@<            �X@������������������������       �2�p@ӽ�?�             s@                          �1@��O���@�           H�@������������������������       ��+��{� @w            �g@������������������������       �:��6��@-           �~@                          �?@�i��@H           ��@                           �?2a�!��@           ��@                          �8@�����^@           `{@������������������������       �z�v�'@�             k@������������������������       �Y!��m@�            �k@                           @a��	@�           �@������������������������       �f�b��		@s           ��@������������������������       �����:@x            �f@                            @/�`^	@F            �^@                           @�˺���@/             V@������������������������       �[���@!             M@������������������������       �[M^u@             >@������������������������       �`;�6G@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        ,@     �r@     ��@      >@     �K@     @~@      V@     ��@     �j@     ��@     �v@     �@@      @     �]@     �r@      1@      3@     �n@     �@@     8�@     �W@     `}@      e@      (@      @      R@     �d@      ,@      0@     @d@      ;@      n@     �R@      k@     �[@       @              7@     �H@      �?       @     �C@      @     �_@      .@     @V@      8@      �?              @      3@      �?       @      :@      @     �Q@      $@      D@      @      �?              1@      >@                      *@              L@      @     �H@      1@              @     �H@      ]@      *@      ,@     �^@      7@     @\@      N@     �_@     �U@      @      @      E@      S@      @       @     @V@      3@     @P@     �D@     �R@     �N@      @              @      D@      @      @      A@      @      H@      3@      J@      9@                     �G@     �`@      @      @     @U@      @     p}@      4@     �o@      M@      @              &@     �B@              �?      6@             �k@      &@     �T@      0@      �?              @      .@                      @             �C@      @      8@      @                      @      6@              �?      1@             �f@      @     �M@      (@      �?              B@     �W@      @       @     �O@      @     `o@      "@     `e@      E@      @               @      4@              �?      (@             �V@      �?      H@       @                      <@     �R@      @      �?     �I@      @      d@       @     �^@      A@      @      "@     @f@     �p@      *@      B@     �m@     �K@     �r@     �]@      r@     �h@      5@      @      d@     �o@      &@      @@     �j@     �H@     `r@     �Z@     0q@      f@      4@      �?      D@     �R@      @      @     �I@      @     �\@      ,@     @W@     �A@      @              9@      B@      @              8@      �?     �O@      �?      K@      $@              �?      .@      C@              @      ;@      @      J@      *@     �C@      9@      @      @      ^@     �f@       @      <@     @d@     �F@     `f@      W@     �f@     �a@      0@      @     @Y@     �b@      @      <@     �`@      D@     �b@     �P@     �c@     ``@      *@       @      3@      @@       @              >@      @      ?@      9@      7@      $@      @       @      2@      (@       @      @      8@      @      @      (@      .@      7@      �?              1@       @               @      $@      @      @       @      (@      5@      �?              ,@      @               @      @      @      @      @       @      *@      �?              @      �?                      @       @              �?      $@       @               @      �?      @       @       @      ,@              �?      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?o�R@�e@�	           ��@       	                    �?��a�U@�            �@                           �?j��b�@%           �}@                            �?-l�qơ@�            �m@������������������������       �W0n���@             J@������������������������       �fc\���@o            @g@                            @��)\�E@�            �m@������������������������       ��y�K�@a            @c@������������������������       � �G��@6            �T@
                          �=@wCH���@�           0�@                           @A�5�n@�           ��@������������������������       ���r�u�@�            pt@������������������������       �&�X� @�            �x@������������������������       �>��_�@             0@                            @_S{u\@�           �@                           �?��f��@�           ��@                            �?0�.��		@Q            ``@������������������������       �*�H�@@            @Z@������������������������       �H��`��@             :@                           @$SN<k�@d           ��@������������������������       �1��(	@&           �@������������������������       �~>�=�#@>            �@                           �?�(3 �	@�           �@                           �?D�h�	@=           �@������������������������       �E��D�	@o            `e@������������������������       �	��y�@�            `u@                           �?Ğýn@�             r@������������������������       ��~�D@             <@������������������������       ���4��@�            `p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     �q@     p�@     �C@      G@     �|@     �W@     ��@     �k@     H�@     �v@     �B@              S@     `b@      @      @     �Y@      0@      |@      B@     `r@     �S@       @             �G@     �Q@      @      @      N@      @     @Z@      9@     @[@     �E@      @              6@      ?@      @      �?      @@      @     �H@      4@     �H@      8@      @              @       @              �?      @       @      ,@      �?      *@       @                      0@      7@      @              ;@       @     �A@      3@      B@      6@      @              9@     �C@               @      <@              L@      @      N@      3@       @              .@      3@              �?      7@              A@      @     �G@      $@       @              $@      4@              �?      @              6@       @      *@      "@                      =@     @S@              @     �E@      (@     pu@      &@      g@      B@      @              =@     @S@              @     �C@      (@     `u@      @     �f@     �@@      �?              1@     �C@              �?      ,@      &@     �a@      @      T@      5@                      (@      C@               @      9@      �?     @i@      @     �Y@      (@      �?                                              @              �?      @       @      @       @      1@      j@     �w@      B@      D@      v@     �S@     ��@     `g@     �@     �q@      =@      "@      a@     �o@      4@      ;@     �n@      L@     @{@     �`@     �v@      i@      .@      @      "@      $@              "@      9@      @      ,@      *@      ;@      *@               @      @      @              "@      6@      @      &@      *@      4@      $@              @      @      @                      @              @              @      @              @     �_@     @n@      4@      2@     �k@     �I@     `z@     �]@     0u@     `g@      .@      @     �R@      ^@      .@       @     �`@     �E@     �`@     @V@      `@     �Z@      *@              J@     �^@      @      $@     @U@       @      r@      >@     `j@     @T@       @       @     @R@     �_@      0@      *@     @[@      6@     ``@     �K@     �b@     �U@      ,@       @      M@     �S@      *@      $@     �T@      0@     �L@      C@     �U@     �I@      ,@      @      ;@      >@      (@      @      >@      @      .@      @      .@      1@      @      @      ?@     �H@      �?      @     �J@      "@      E@      ?@     �Q@      A@      &@              .@      H@      @      @      :@      @     �R@      1@     �O@     �A@                      @      @              �?              @      �?      @              @                      &@     �D@      @       @      :@      @     @R@      $@     �O@      >@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJs�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@H6�u@�	           ��@       	                   �1@�C��4@           t�@                           @(�2df�@�           ��@                           @�D/��Q@�            �o@������������������������       �09e��@�             n@������������������������       �������@	             .@                           @�	}��
 @�            �u@������������������������       ��A��_�?�            �p@������������������������       ��2J�D�@5             U@
                          �5@�Ѭ��@�           x�@                            �?�����@�           �@������������������������       �Mb���3@�            @v@������������������������       ��"c 6@�           x�@                            �?Q�G�}@�            �u@������������������������       ���R=�@:            �Y@������������������������       �#Xw��2@�            �n@                           @���)�@�           <�@                          �;@�N��n�	@Y           ��@                           �?I/s��@�           0�@������������������������       ������@(           �|@������������������������       �Jd�z@f            `c@                            �?^����	@�            �r@������������������������       ��m�1�	@e            `b@������������������������       �z��~�@f             c@                           @*]̝l@2           �@                           @Ϟ��˴@            {@������������������������       ���F�T�@�             p@������������������������       �4Ƞ���@g            @f@                          �:@Ş�'ʺ@-            �R@������������������������       �?h�i@             J@������������������������       �S���% @             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@      r@     ��@      ?@      P@     �@      U@     �@      j@     ��@     �v@      A@      *@     �c@     �v@      3@     �@@     �q@      @@     P�@     �Y@     p@     �g@      *@              4@     �U@       @      @     �H@       @      p@      3@      `@      A@                      0@      E@       @              >@       @     �T@      1@      E@      5@                      ,@      D@       @              8@             �T@      0@      E@      4@                       @       @                      @       @      �?      �?              �?                      @     �F@              @      3@             �e@       @     �U@      *@                      @      <@                      $@             @a@      �?     @R@      &@                              1@              @      "@             �A@      �?      ,@       @              *@     @a@     0q@      1@      ;@     �m@      >@     P�@      U@     `w@     �c@      *@      &@      W@      k@      .@      3@      h@      :@     @{@     �P@     �s@     �`@      *@              5@     �D@              �?     �I@      @     �Y@      .@     �V@      ;@      @      &@     �Q@     �e@      .@      2@     �a@      7@     �t@      J@     @l@      [@      "@       @      G@     �M@       @       @      F@      @     �U@      1@      M@      6@               @      8@      ,@      �?      @      $@              <@      @      @       @                      6@     �F@      �?      @      A@      @      M@      $@      K@      ,@              "@     @`@     @f@      (@      ?@     �k@      J@     `n@     �Z@      o@     @e@      5@      "@     �W@     �]@      $@      2@     �d@     �F@      ]@     �S@     @]@      _@      4@              L@     �R@      @      $@     �]@      <@     �X@     �J@     �V@      P@      1@             �D@      M@      @       @      Z@      2@      O@      G@      O@     �C@      0@              .@      0@               @      .@      $@      B@      @      <@      9@      �?      "@      C@      F@      @       @     �F@      1@      2@      :@      ;@      N@      @      @      "@      5@       @      @      .@      &@      @      1@      2@     �A@       @      @      =@      7@      @      @      >@      @      (@      "@      "@      9@      �?              B@      N@       @      *@      M@      @     �_@      ;@     �`@      G@      �?              6@      F@       @      *@     �H@      @     @\@      2@     @_@     �E@                      &@      =@              @      9@             �Q@      @     �U@      6@                      &@      .@       @      "@      8@      @      E@      &@      C@      5@                      ,@      0@                      "@       @      ,@      "@      @      @      �?              @      .@                       @       @      *@      "@      @       @      �?              $@      �?                      @              �?              @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���F&]@�	           ��@       	                     @O��	�I@�           �@                          �0@��9�[�@N           $�@                            �?�As�}��?b            �d@������������������������       �z���  @E            @^@������������������������       ��0��^�?             G@                           �?��s�m�@�           ��@������������������������       ���xd@^           ��@������������������������       �Dqh�*@�           X�@
                          �2@J�5�@2           �@                           @lJ9�&�@�            �t@������������������������       ��m�
g@�             l@������������������������       ��3��	�?:            �Z@                           �?����Q@v            `f@������������������������       �+�Z�@J            �Z@������������������������       ��psl�@,            @R@                          �<@/��P�@           �@                           �?��8
�X@P           d�@                           �?�����	@�           h�@������������������������       ��5�B��	@�            Ps@������������������������       �!8��
	@!           �}@                           �?��##��@g           `�@������������������������       ��u^S:@�            0q@������������������������       �u�R��@�           ȅ@                          �?@��X�[�@�            �r@                            @�Ǜ��@�            @i@������������������������       �^���K@Y            �a@������������������������       �lކ��@*             N@                          @A@_6��m]	@?            �W@������������������������       �e_r~@4            �S@������������������������       �Ii��G@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     0s@      �@      =@     �M@     �z@      S@     @�@     �l@     �@      v@      A@       @     �X@     �q@      @      2@     @f@      *@     ��@     @U@      x@     �a@      "@              R@     `k@      @       @      `@      @     �~@     �P@     �p@      T@      @              �?      E@                      $@              S@              ;@      &@                      �?      =@                      @              L@              1@      &@                              *@                      @              4@              $@                             �Q@      f@      @       @     �]@      @     z@     �P@      n@     @Q@      @              <@      S@       @      @      M@             @i@     �E@     @W@      =@      �?             �E@     @Y@      @      @     �N@      @     �j@      8@     `b@      D@      @       @      :@     �P@       @      $@     �H@      @     �a@      2@     �]@      N@       @       @      .@     �C@      �?      @      C@             @Y@      "@     �T@      C@               @      *@      @@      �?      @      :@             �J@      "@     �H@      A@                       @      @                      (@              H@             �@@      @              @      &@      ;@      �?      @      &@      @      E@      "@     �B@      6@       @      @      $@      $@               @      @      @      .@      "@      =@      ,@       @              �?      1@      �?       @      @       @      ;@               @       @              &@      j@     0r@      6@     �D@     @o@     �O@     �v@      b@     �y@     �j@      9@      $@     �f@     p@      2@      <@     �i@      J@     �u@      \@     �v@     �c@      7@      $@     @Z@      ^@      .@      *@     @]@      8@      V@      P@      `@     @T@      0@      @     �G@      J@      $@      @     �D@      "@      G@      2@     �@@      B@      @      @      M@      Q@      @      @      S@      .@      E@      G@     �W@     �F@      $@             �R@      a@      @      .@     @V@      <@     p@      H@     �m@     @S@      @              0@      B@      �?              4@      @     @\@      @     @R@      $@                     �M@     @Y@       @      .@     @Q@      9@      b@     �F@     `d@     �P@      @      �?      =@      A@      @      *@      F@      &@      3@     �@@     �I@      L@       @              0@      7@              "@      <@      "@      .@      9@      >@     �G@                      @      $@              @      5@      @      &@      2@      6@     �C@                      "@      *@               @      @       @      @      @       @       @              �?      *@      &@      @      @      0@       @      @       @      5@      "@       @              (@      @       @      @      *@      �?      @       @      3@       @       @      �?      �?      @       @              @      �?                       @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�.�5h@�	           ��@       	                    �?[ְj	@�           h�@                           �?oY0&�@~           �@                          �2@�*�@�            q@������������������������       �������@*            @S@������������������������       �B���J@v            �h@                           �?��
X�@�             u@������������������������       ��!�E�@K             \@������������������������       ���[��4@�             l@
                            �?;�+��	@t           ȏ@                          �7@��!�C�	@�             r@������������������������       � `��S�@g             e@������������������������       ��@pD�)	@H             ^@                          �;@"}����	@�           Ȇ@������������������������       �ä���	@t           ��@������������������������       ���9d�@Q            �`@                          �3@����@�           ޡ@                           �?	���j@j           �@                           �?��E�K�?�            �w@������������������������       �?�G�e��?�            �h@������������������������       ��
5#:�?l            �f@                           @Y>(&�@~           8�@������������������������       ��\���@�            �o@������������������������       �����@�            �v@                           �?'���X`@;           0�@                          �=@��S��:@�            `x@������������������������       �ͳ0tuy@�            w@������������������������       ��X�x@             5@                          �<@��)&7I@L           0�@������������������������       ��r�"@           ��@������������������������       �ǣ-��@:            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �p@     ��@      C@      N@     P|@     �U@     �@     @l@     p�@     pv@      >@      3@      b@     �o@      ?@      D@     `o@      H@     @l@     �`@     �o@     �i@      5@      @     �A@     @Y@      @      &@     �W@      $@     �^@      G@      Z@     �Q@      @      @      3@      F@      @      �?     �K@      @     �O@      0@     �B@      5@      @      @      @      *@                      *@      �?      A@              @      @              �?      .@      ?@      @      �?      E@      @      =@      0@      @@      1@      @              0@     �L@      �?      $@     �C@      @     �M@      >@     �P@      I@       @              @      3@                      ,@              9@      @      >@      ,@                      "@      C@      �?      $@      9@      @      A@      ;@     �B@      B@       @      .@     @[@      c@      ;@      =@     �c@      C@      Z@     �U@     �b@     �`@      ,@      �?     �E@     �D@      @      $@      D@      &@      :@     �A@     �H@      5@      @              7@      5@               @     �@@       @      4@      ,@      ?@      1@      @      �?      4@      4@      @       @      @      "@      @      5@      2@      @              ,@     �P@      \@      5@      3@     @]@      ;@     �S@      J@      Y@     �\@      "@      "@     �I@      W@      1@      $@     @Y@      6@     �R@      G@     �U@     @S@      "@      @      .@      4@      @      "@      0@      @      @      @      *@     �B@                      ^@      t@      @      4@     @i@     �C@     ؇@     @W@     ��@      c@      "@              ?@     @^@      @      @     �N@      �?     �y@      D@     �p@     �G@       @              .@      =@                      @             `h@      "@     @\@      $@       @              @      *@                      @             @\@      @     �H@       @                      "@      0@                      @             �T@      @      P@       @       @              0@      W@      @      @      K@      �?     @k@      ?@     �c@     �B@                      "@      I@               @      5@      �?     �T@      <@     �C@      4@                      @      E@      @      @     �@@             �`@      @     �]@      1@                     @V@     �h@      @      ,@     �a@      C@     �u@     �J@     0r@     �Z@      @              *@     �P@                     �@@      &@     �b@       @      V@      5@                      *@     @P@                      =@       @     @b@      @     �U@      2@                               @                      @      @      @      @      �?      @                      S@     �`@      @      ,@      [@      ;@      i@     �F@     `i@     @U@      @              Q@     �^@      @      ,@     @V@      7@     �g@     �E@      h@      R@      @               @      $@      �?              3@      @      &@       @      $@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-�RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��
Ռ@@�	           ��@       	                    @�����`@           4�@                          �<@y���B@�           ��@                           �?�^Lp�@q           ؁@������������������������       ��#�K5@           �y@������������������������       �l����@l             d@                           �?�l�l�m@,             Q@������������������������       ���=h�@
             3@������������������������       ����3�t@"            �H@
                          �2@�9HC&@y           p�@                            �?qlq��?�            @n@������������������������       �`m����?M             _@������������������������       �}�K��?G            �]@                            @pe�M0@�            �u@������������������������       ��'��o@�            @r@������������������������       �y(�[�P�?"             L@                           @r}^�B,@�           ��@                          @A@�I��lq	@�           @�@                          �3@9y� H	@�           �@������������������������       ��ξ���@           �{@������������������������       �3�:�܇	@�           �@������������������������       �jg���@	             .@                          �7@yZ4�7�@�           ��@                          �1@����@           x�@������������������������       �ͯ�sO @w            �g@������������������������       ���QԞ@�           ��@                           @�dƬiO@�            �q@������������������������       ����W�@�            �l@������������������������       �`���T@$            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        .@     �r@     ��@      5@      K@     �~@     @T@     �@      j@     ��@     �w@     �@@              Q@     �c@       @      &@     �]@      "@     �{@      C@      r@     @V@      @             �I@     �T@       @       @      S@      @     �b@      <@      e@     �P@      @             �G@     �R@       @      @     �O@      @     �a@      5@     �d@     �F@      @             �A@     @P@       @      @      H@      @     �U@      3@     @[@      B@      @              (@      $@              �?      .@      @      K@       @     �K@      "@                      @      @              @      *@              @      @      @      5@      �?               @      @                       @              @                      @                       @       @              @      &@               @      @      @      0@      �?              1@     �R@              @     �E@      @     pr@      $@      ^@      7@      �?               @      7@               @      .@             �b@      @      @@      @      �?              @      &@               @      "@              T@              (@      @                       @      (@                      @             �Q@      @      4@              �?              "@      J@              �?      <@      @      b@      @      V@      3@                      "@      H@                      8@      @      \@      @     �R@      1@                              @              �?      @              @@              *@       @              .@     �l@      x@      3@     �E@     pw@      R@     0�@     @e@     �@     0r@      <@      .@      c@     �l@      0@      C@     �o@     �P@      i@     ``@     @l@      i@      7@      $@     �b@     �l@      *@      C@     �o@     @P@      i@     @`@     @l@     �h@      7@      @      =@     @P@      @      @     @P@       @     �V@      E@     @Q@     �N@      �?      @     �^@     �d@      $@      @@     �g@     �L@     @[@      V@     �c@      a@      6@      @       @              @                      �?              �?              @                     �S@     `c@      @      @     �^@      @     �u@     �C@     `q@     �V@      @              H@     �`@      @      @      O@      @     �r@      4@     `j@     �O@       @              @      =@                      @             �T@      @     �K@      "@                      E@     �Z@      @      @      M@      @     �j@      1@     �c@      K@       @              >@      4@               @      N@       @      K@      3@     �P@      <@      @              2@      (@               @      J@      �?     �E@      (@      P@      8@                      (@       @                       @      �?      &@      @      @      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�J>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �2@�_�kr�@�	           ��@       	                    @`%b�G@�           Ȑ@                           @]�%$�@            �@                            @Q+}���@�            �x@������������������������       ��D�Q� @�            �m@������������������������       �>u(�w@f            �c@                          �1@`F�*�� @           �}@������������������������       �.��P�s�?�            �r@������������������������       ����i�)@m            �e@
                           @X��wh@�            @j@                          �0@d7qt}@}            �h@������������������������       ��C�3���?              K@������������������������       �����v@]             b@������������������������       ��tc��@             &@                           �?���C^@           .�@                           �?��i�}@�           �@                            �?c��R�@�            `t@������������������������       �野�x@v            @f@������������������������       ���*�f@\            �b@                           @�w�E5t@*           �}@������������������������       �����"@S            �_@������������������������       ��1��f=@�            �u@                          �9@��/�	@           П@                           @�YBr{@�            �@������������������������       �<�b�w1@v           ��@������������������������       ��p�Vd�@G           �~@                           �?8��x��	@a           ��@������������������������       ��|�.u
@�            �r@������������������������       �>��XY>@�            Pp@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        6@     �r@     ��@     �D@      L@     �{@      V@      �@      j@     ��@      y@      ?@      @     �J@     �_@       @      $@     �W@       @     @z@     �D@     �l@     �T@       @             �A@     �X@       @       @     �S@      @      u@      >@     `j@      M@      �?              5@      F@      �?      @      J@      @     @[@      7@     @U@     �G@                      $@      2@                      A@             �S@      0@      J@      <@                      &@      :@      �?      @      2@      @      ?@      @     �@@      3@                      ,@      K@      �?      @      ;@      �?     `l@      @     �_@      &@      �?              "@      ?@                      1@             �b@             @T@       @      �?              @      7@      �?      @      $@      �?      S@      @     �F@      @              @      2@      =@               @      .@       @      U@      &@      4@      8@      �?      @      2@      <@               @      &@             �T@      &@      2@      8@                      �?      *@                      @              =@              @      @              @      1@      .@               @      @              K@      &@      ,@      5@                              �?                      @       @      �?               @              �?      2@     �n@     py@     �C@      G@     v@      T@     ��@      e@     ��@      t@      =@              S@     �_@       @       @     @Q@      "@      k@      A@      i@      P@      @             �I@     �L@       @      �?     �@@      �?     �G@      7@     @Q@      D@       @              7@      >@       @      �?      (@              <@      "@     �F@      :@       @              <@      ;@                      5@      �?      3@      ,@      8@      ,@                      9@     �Q@              �?      B@       @     @e@      &@     ``@      8@      �?              (@      .@                      &@      @     �B@      "@      @@      @      �?              *@     �K@              �?      9@      @     �`@       @     �X@      3@              2@     @e@     �q@     �B@      F@     �q@     �Q@     0v@     �`@     �v@      p@      :@       @     �]@     �j@      8@      =@     �i@     �F@     �r@     @U@     pq@     �b@      0@      @     @P@     �^@      2@      5@      b@     �@@     �k@     �C@     @h@     �Y@      &@       @     �J@     �V@      @       @      N@      (@     �S@      G@     @U@     �G@      @      $@      J@     �P@      *@      .@      T@      :@     �J@     �H@     �T@     �Z@      $@      $@      =@      A@      "@      @     �E@      6@      *@      :@      @@     �Q@      $@              7@     �@@      @      $@     �B@      @      D@      7@      I@     �B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�p�@�	           ��@       	                    @T%H��@�           ��@                           �?ҩe�@<           ��@                           �?�|��R�@�           Ȃ@������������������������       �$^����@�             n@������������������������       ���#��x@�            �v@                          �3@�S�l�z@�            �q@������������������������       ��Eo�@�            `m@������������������������       ���zЕ@%             J@
                           �?ל��+@\           `�@                          �0@��ه���?�            @v@������������������������       �%�X��� @              L@������������������������       �.��.���?�            �r@                          �1@	�P5�@t           @�@������������������������       �#�}2�9�?�            �h@������������������������       ��`��@�            @x@                           @��xK0@2           J�@                           �?�����@F           H�@                          �<@ulEb�@�            w@������������������������       �2Q�U|@�            �r@������������������������       �{�@*             Q@                           @\9���&	@W           �@������������������������       �'�6v¹@           @�@������������������������       ���� 
@K            @^@                          �8@�{7n�@�           ��@                           @��[@)           �}@������������������������       �Z����@B            �X@������������������������       ��L��@�            `w@                           @��"&��@�            �s@������������������������       �p�@'�@�            �r@������������������������       ��/�Q�@	             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     P�@     �A@     �E@     �{@      S@     ��@     �i@     ��@      t@      :@       @     �Y@     �n@      (@      *@     `e@      *@     8�@      V@     �x@     �_@      @       @      O@     @`@      @      @      ^@       @     @l@     �Q@     �d@     �T@      @       @     �H@     @T@      @       @     �V@      @     �a@      F@     �Y@     �P@      @       @      3@      G@      @             �B@      @     �P@      0@      =@      1@      �?      @      >@     �A@      �?       @     �J@      @      S@      <@     @R@      I@      @              *@     �H@       @      @      >@      �?      U@      :@      O@      0@                      *@      B@              �?      2@      �?     �R@      7@      L@      *@                              *@       @      @      (@              $@      @      @      @                     �D@      ]@      @      @     �I@      @     Pz@      2@      m@     �E@      �?              "@     �C@               @      .@             �h@      @     @S@      "@      �?                      (@                      @              5@              *@      @                      "@      ;@               @      "@             @f@      @      P@      @      �?              @@     @S@      @      @      B@      @     �k@      *@     `c@      A@                      @      8@              @      @             �X@             �M@      @                      =@     �J@      @       @      @@      @      _@      *@      X@      =@              &@      j@     @s@      7@      >@     �p@     �O@     �y@     @]@     �z@     @h@      5@       @     �d@     �g@      .@      7@      i@     �J@     �f@     @V@      l@     �`@      .@      �?     �G@     �E@      @      $@     �H@       @     �T@      2@     @T@      ;@      @      �?     �E@      ?@      @       @     �B@       @      T@      "@     �Q@      ,@       @              @      (@               @      (@               @      "@      &@      *@      @      @     �]@     `b@      &@      *@      c@     �I@     �X@     �Q@     �a@     �Z@      $@      @     @Z@      `@      @      (@     �a@     �F@      T@      J@     �`@     @W@      @      �?      ,@      2@      @      �?      (@      @      3@      3@       @      *@      @      @     �E@     �]@       @      @      Q@      $@      m@      <@     `i@     �N@      @      @      >@     �U@      @      �?     �F@      @     �a@      $@      \@      <@      @      @      �?      5@       @               @      @      =@      �?      6@      @      @              =@     �P@       @      �?     �B@       @     @\@      "@     �V@      6@      @              *@      ?@      @      @      7@      @     �V@      2@     �V@     �@@                      "@      >@      @      @      3@      @     �V@      1@      V@     �@@                      @      �?                      @      �?              �?      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJpF/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�b��@�	           ��@       	                    �?}:y�5�@u           B�@                          �;@H��-	@�           ��@                           @Xx��@V           ��@������������������������       �aU��l@G           X�@������������������������       �2�&��@             :@                           �?�a��
@�             o@������������������������       ��"&C��@*            @Q@������������������������       �o`��.
@y            �f@
                           �?l_�k��@|           ��@                          �1@�����>@�            �p@������������������������       �k\��v @            �C@������������������������       ���9��@�            `l@                           �?�bP�A@�            �v@������������������������       ��pF@5            �U@������������������������       �6����@�            �q@                           �?E^��Z�@L           ��@                           @�3��'��?t           ��@                          �4@O�%��?�            �s@������������������������       ��Ʉ1-m�?�            �i@������������������������       �e�!.@C             [@                            @O	j��a @�            �o@������������������������       ���"6l[ @�            �g@������������������������       �@��@|��?%             O@                          �1@q��.@�           ȑ@                           �?��	����?�             i@������������������������       �[��`mq@@            @W@������������������������       ��}Eٟ1�?F            �Z@                           @a����@R           P�@������������������������       �j^��@�           p�@������������������������       ��;�i�\@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     @q@     h�@      @@      K@      |@      R@     `�@     �k@     �@     �s@     �A@      4@     `j@     �t@      6@      C@     ps@     �L@     �x@      f@     �x@     �k@      :@      4@     `d@     `m@      4@      ;@     `m@      G@     �l@      `@     0q@     �e@      8@      *@     �`@     @i@      (@      2@     @k@      >@     �i@     �[@     �n@     @]@      5@      "@     ``@     @i@      (@      2@     @j@      <@     �i@     �[@     �n@     @]@      .@      @      @                               @       @      �?      �?                      @      @      <@     �@@       @      "@      1@      0@      7@      1@      ?@     �L@      @       @       @      @      �?       @      @      @      "@              ,@      1@              @      4@      =@      @      @      &@      $@      ,@      1@      1@      D@      @              H@     �X@       @      &@      S@      &@     �d@      H@     @^@      H@       @              2@      =@       @      @      B@      @      Q@      4@     �K@      9@      �?              �?      @                       @              3@      @      @                              1@      7@       @      @      A@      @     �H@      0@      H@      9@      �?              >@     �Q@              @      D@      @     �X@      <@     �P@      7@      �?              @      @                      @              @@      @      =@       @      �?              8@     �O@              @      A@      @     �P@      9@     �B@      5@                     @P@     �k@      $@      0@      a@      .@     `�@      G@     P{@     �W@      "@              (@     �M@      �?      @      8@      @     @s@      *@      `@      (@      �?               @      ?@                      ,@       @      g@      "@     �L@      @                      @      2@                      @             �a@              @@      @                      @      *@                      @       @      F@      "@      9@      @                      @      <@      �?      @      $@      �?     �^@      @      R@      @      �?               @      ;@      �?      �?      $@      �?     @X@      @      F@      @      �?               @      �?              @                      :@              <@       @                     �J@     �d@      "@      (@     @\@      (@     �u@     �@@     @s@     �T@       @              @      >@               @      @             @W@      �?     �L@      @                      @      3@               @      @              E@      �?      2@      @                       @      &@                       @             �I@             �C@       @                      H@     �`@      "@      $@      [@      (@     `o@      @@     `o@     �R@       @              :@     �V@      @      @     @Q@      @     @j@      4@     �e@     �D@      @              6@     �E@      @      @     �C@      @     �D@      (@      S@      A@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ/��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�虀!@�	           ��@       	                    �?zxd�u�@           ԓ@                            @�^*1�@B           �@                           �?�Ƽ�H@�            �r@������������������������       �0f�K�v@O            �_@������������������������       ��?Y`�0@n             f@                           �?�~����@�            �i@������������������������       ����F�.@*             R@������������������������       �I�f�88@[            �`@
                          �>@����@�           ��@                           @,Xʺ}@�           �@������������������������       ��m�I�. @W           ��@������������������������       ����Lq@t            �h@                          @@@�\{�/@             5@������������������������       �E�2�� @             (@������������������������       ���!zȓ@             "@                          �5@��|�A
@�           ��@                            @���9y$@�           l�@                           �?�����W@�           ؐ@������������������������       �����@�             n@������������������������       �/C�H�@�           0�@                          �1@+Gc�0@�            Pv@������������������������       �z�o�@:            @X@������������������������       ��V>kER@�            @p@                           @�]"Dr	@           �@                          �:@2�S���	@�           ��@������������������������       �Z� 1��	@=           �@������������������������       ������k	@�            �q@                          �<@��c AA@           `z@������������������������       �����Ӫ@�            `v@������������������������       ��u��`�@)             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@      �@      2@     �Q@     p{@     �T@     ��@      j@     8�@      v@     �@@      @     �V@     �e@       @      .@      Z@       @      }@      @@     �q@     �T@      @      @      L@      U@       @      "@      O@       @      \@      6@     @[@      F@      @      @      B@     �C@      �?       @     �E@       @     �N@      *@     �P@      ?@      @      @      1@      1@      �?       @      (@       @      =@      "@      .@      2@      �?              3@      6@                      ?@              @@      @      J@      *@      @              4@     �F@      �?      @      3@             �I@      "@      E@      *@                      @      4@                       @              9@      �?      2@       @                      0@      9@      �?      @      1@              :@       @      8@      &@                     �A@     @V@              @      E@      @      v@      $@      f@      C@       @             �A@     �U@              @      B@      @     �u@      @      f@      A@       @              9@     @P@              �?      3@      @     Pq@      @     �_@      4@                      $@      6@              @      1@              R@      @      I@      ,@       @                       @                      @      �?      @      @              @                               @                      @               @      �?               @                                                      �?      �?      @       @               @              *@     �j@     0u@      0@     �K@     �t@     �R@     ��@      f@     H�@      q@      :@      @     �Q@     `i@      @      2@     @e@      :@     z@     @Q@     pt@      ]@      $@       @      G@      d@      �?      &@     �]@      *@     �t@     �I@     p@     �T@      @       @      <@      <@              @     �D@      @     �B@      6@      A@      A@      @              2@     �`@      �?      @     @S@       @     `r@      =@     �k@     �H@      �?       @      9@     �E@      @      @      J@      *@     �U@      2@     �Q@     �@@      @              &@      (@      �?      �?      @             �A@      @      0@      &@               @      ,@      ?@       @      @      H@      *@     �I@      (@      K@      6@      @      "@     �a@      a@      (@     �B@     �d@      H@     `g@      [@     @h@     �c@      0@      "@     �Y@     @W@      "@      8@     �[@     �D@     @T@     �U@     @Z@     �[@      ,@      @     �Q@     �Q@      @      2@     @R@      8@     �M@     �K@      S@     �D@      $@      @      ?@      6@      @      @      C@      1@      6@      @@      =@     �Q@      @             �C@     �E@      @      *@      K@      @     �Z@      5@     @V@     �F@       @              =@      C@       @       @     �B@      @     �Z@      4@     @S@      @@       @              $@      @      �?      @      1@                      �?      (@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ/�m@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @YuRy�H@�	           ��@       	                    �?/�F��@�           ��@                          �;@�H�z�@�           �@                            �?���2F@i           @�@������������������������       �ޝ�<�u@x            `i@������������������������       �	�o�z@�            �w@                          �<@'�{�B@7            �V@������������������������       �V@���@             *@������������������������       ��K���@/            �S@
                           �?�c7�%5	@�           ��@                          �9@x!p�37	@M            �\@������������������������       �Ne�S@5            @S@������������������������       �����@            �B@                           @�76	@�           ܖ@������������������������       �Pý��@�           `�@������������������������       ���Us<q	@           X�@                           @=��$qL@           ��@                           @��v@�           ��@                           �?��Щ��@�           ��@������������������������       ��W�N\�@�             {@������������������������       �-{�7C@�           ��@                           @�I>U��@B           �@������������������������       �d�>H@�            �p@������������������������       �p\���@�            `n@                           @� kǝX@             9@������������������������       �-�Nk�t@             .@������������������������       ������@	             $@�t�bh�h5h8K ��h:��R�(KKKK��h��B 
        .@     `t@     h�@      ;@      F@      }@     �W@     `�@     �m@     p�@     0u@      6@      .@     `m@     �u@      5@      ;@     �t@     �R@     0x@      h@     �w@     �k@      3@      �?     @Q@     �W@       @      @     @X@      @     �e@      8@      c@      I@      @             �J@     �U@       @       @     @T@       @      d@      1@      a@     �D@      @              (@      A@                      9@      �?      J@      @      M@      .@       @             �D@      J@       @       @      L@      �?     @[@      *@     �S@      :@      �?      �?      0@      "@              @      0@      @      &@      @      0@      "@              �?      @                                      @      @               @                              (@      "@              @      0@               @      @      ,@      "@              ,@     �d@     �o@      3@      6@      m@     @Q@     �j@      e@     `l@     �e@      0@      @      1@      $@              @      3@      @      @      5@      2@      @       @      �?      $@      @              @      1@      @      @      &@      *@      @              @      @      @                       @      �?              $@      @      �?       @      "@     �b@     �n@      3@      2@     �j@     @P@      j@     `b@      j@     �d@      ,@       @     �L@     @Z@      @       @     @X@      @@      Y@      A@     �Y@      T@       @      @      W@     �a@      (@      0@     @]@     �@@      [@     @\@     �Z@     �U@      (@             �V@     �i@      @      1@     �`@      4@     H�@     �G@     0{@      ]@      @             �T@     �i@      @      0@     ``@      0@     @�@      F@      {@      ]@      @             �L@     `b@      �?      @      U@      &@     �{@      5@     �r@     �N@       @              5@      N@                      7@      &@     �h@      @     �Y@      *@                      B@     �U@      �?      @     �N@             �n@      .@     @h@      H@       @              :@     �M@      @      *@     �G@      @     �a@      7@      a@     �K@      �?              @      >@       @      "@      2@      @      V@      3@     �P@      8@                      4@      =@       @      @      =@      �?     �J@      @     @Q@      ?@      �?               @      �?      �?      �?      @      @      �?      @      @                              @              �?              @      @              @                                      @      �?              �?              �?      �?              @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ<+ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�.~~�B@�	           ��@       	                    �?��K@�@u           ֠@                           �?��4m@�           `�@                          �2@�^�߷�@�            pp@������������������������       ���$�o$@P            �_@������������������������       ���6I�@[             a@                           �?�\�q	@<           P~@������������������������       ���K!�@e             e@������������������������       ��M�QE�@�            �s@
                           �?����Y�@�           ��@                          �0@�G�%wG @7           p~@������������������������       �08�^��?%             P@������������������������       ��E�!��?           pz@                            �?9Ɲ8��@W           ��@������������������������       ��(z	�H@�             k@������������������������       �FP�ğ�@�           ��@                           �?T�0ς�@V           x�@                            �?g6�J@�           ��@                          �9@�BS�	@z            �g@������������������������       �+�ᛕ�@M            @^@������������������������       ����d�@-            �Q@                           @�)4\O\@L           ��@������������������������       ���75�a@�            0s@������������������������       ��8П�L@�            @l@                            �?g-w]�@�           (�@                           @���eJ	@\           �@������������������������       ��F����	@�            w@������������������������       ���D�Du@m             f@                          �<@X�;g�@4           �~@������������������������       ���? @�            �x@������������������������       �ngX�D@;            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     pt@     ȁ@      =@      M@     �y@     �Q@     ��@     �k@     (�@     pv@     �@@      "@     �[@     @s@      @      <@     �k@      9@     ��@     �U@      @     `c@      .@      "@      N@     �W@       @      ,@     �[@      (@     `b@     �L@     `c@     @S@      $@              3@      A@      �?      �?      @@              T@      (@     �P@      0@      �?              @      .@                      :@             �E@      @      ;@      @                      .@      3@      �?      �?      @             �B@      @      D@      $@      �?      "@     �D@      N@      �?      *@     �S@      (@     �P@     �F@      V@     �N@      "@      @      (@      =@      �?      @      9@      @      8@      (@      8@      :@              @      =@      ?@              "@      K@      @     �E@     �@@      P@     �A@      "@             �I@     �j@      @      ,@      \@      *@      �@      >@     Pu@     �S@      @              3@     @R@              @      7@             �o@      @      X@      *@      �?                      8@                      @              8@               @       @                      3@     �H@              @      1@             �l@      @      V@      &@      �?              @@     �a@      @      &@     @V@      *@     0r@      8@     �n@     @P@      @              @      B@                      0@       @     �U@      &@     �E@      1@                      :@     @Z@      @      &@     @R@      &@     �i@      *@     @i@      H@      @      @      k@     Pp@      6@      >@      h@      G@      t@     �`@     Ps@     �i@      2@             @W@     @^@      &@      .@     �R@      1@     `b@     �F@      \@     @T@      @              1@      =@               @      ?@      @      J@      0@      8@      *@      @              *@      ,@                      8@              C@      $@       @      &@      @              @      .@               @      @      @      ,@      @      0@       @                      S@      W@      &@      *@      F@      *@     �W@      =@      V@      Q@      @             �M@     �K@      $@      @      9@      "@      6@      2@      H@      J@      @              1@     �B@      �?      @      3@      @     @R@      &@      D@      0@      �?      @     �^@     �a@      &@      .@     @]@      =@     �e@     @V@     �h@     �^@      &@      @     @R@     @Q@       @      (@      M@      1@     �P@     �J@      [@     �P@       @      @     �L@      G@      @      (@      D@      ,@      9@     �C@     �P@      I@       @              0@      7@       @              2@      @      E@      ,@     �D@      1@              �?      I@     �Q@      @      @     �M@      (@     �Z@      B@     @V@      L@      @      �?      A@     �N@       @       @     �E@      "@     �W@      =@      U@     �A@      @              0@      $@      �?      �?      0@      @      &@      @      @      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�3,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @8��1�S@�	           ��@                          �2@|,�%�@w            �@                           @U��;W6@*           @                           �?ˢ x��@           `}@������������������������       �Y���@�            Ps@������������������������       �7����a@a             d@������������������������       ��q7t`�@             ;@                           �?�k�h	@M           |�@	       
                    �?��p[pd@"           �z@������������������������       ��2���@w             f@������������������������       ��]�;ܞ@�            `o@                          �@@y�B�ޜ	@+           ̓@������������������������       ��:}߮�	@           \�@������������������������       �9	"�q@             <@                          �6@_ ���@$           �@                           �?��N#�{@�           ��@                          �2@��t�@�           (�@������������������������       ��js_� @�            �r@������������������������       ���v�_@�            �u@                          �1@v#$�(@Z           P�@������������������������       �Kw��k��?c             e@������������������������       � !�◐@�             x@                           @�ʭ�k@:           P�@                           @M�[	 @�            �t@������������������������       �phJ2��@�             l@������������������������       ���	4��@?            �Z@                           @r��0@r            �g@������������������������       �	<�>Y�@7             V@������������������������       ��-b�@@;            �Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     �r@     0�@      A@     �O@     �{@      T@     ��@     �j@     �@     �v@      8@      1@     `l@     @s@      8@     �H@     �r@      Q@     pw@     @f@     0w@     @p@      3@       @      C@      P@      @      �?      L@      @     �a@      A@     �X@      J@               @     �B@     �N@      @      �?     �G@      �?     �a@      @@      W@     �I@               @      =@     �C@      @      �?     �B@      �?     @S@      3@      O@      C@                       @      6@                      $@             @P@      *@      >@      *@                      �?      @                      "@      @      �?       @      @      �?              .@     �g@     �n@      4@      H@      n@     �O@      m@      b@     q@      j@      3@              A@     �O@      @      $@     @P@      .@      S@      >@      T@      G@       @              ,@      4@      @      �?      =@      @      ?@      0@      D@      2@      �?              4@     �E@      @      "@      B@      &@     �F@      ,@      D@      <@      �?      .@     `c@     �f@      *@      C@     �e@      H@     �c@     �\@      h@     @d@      1@      (@      c@     @f@      *@      B@      e@      F@     �c@     �\@      h@     `c@      1@      @       @      @               @      @      @                              @               @      R@     @n@      $@      ,@     �b@      (@     �@     �A@     �|@     �Z@      @              ?@     `e@      @      (@     @U@      @     �}@      1@     �t@     �N@      @              *@      R@      @      $@     �P@      @     p@      (@     �d@      D@                      @     �D@      �?      @      2@              a@      @     �T@      "@                      "@      ?@      @      @      H@      @     @^@       @      U@      ?@                      2@     �X@               @      3@              k@      @      e@      5@      @                      9@                      @             �O@       @     �P@      @       @              2@     �R@               @      (@             @c@      @     �Y@      2@       @       @     �D@     �Q@      @       @     �P@      "@     �`@      2@      `@     �F@      �?       @      =@     �F@                     �D@      @      W@      @     �U@      9@      �?       @      *@      =@                      ;@      @     @R@       @     �O@      &@                      0@      0@                      ,@              3@      @      7@      ,@      �?              (@      :@      @       @      9@      @     �E@      *@      E@      4@                              2@      @      �?       @      �?      >@      $@      3@      @                      (@       @              �?      7@      @      *@      @      7@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�0xBhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @a���ς@|	           ��@       	                    �?��U�@c           0�@                           �?1��_@�           ��@                          �8@E�@/           }@������������������������       ��}=E@�            @u@������������������������       �)[����@R            @_@                            �?��D�p@v            �e@������������������������       ��;�wQ� @%             J@������������������������       ����a�/@Q            �^@
                           @��GOy	@�           d�@                           �?9MqS	@K           p�@������������������������       �hw8]b@�            �v@������������������������       ���r�B�	@g           ��@                            �?Sn��	@s            �g@������������������������       ��~��V/@(             O@������������������������       ���rq�@K            �_@                          �4@=�9R�}@           Ě@                          �1@�gk@*           ��@                           @�:���?�            �v@������������������������       ��I�~B�?�             j@������������������������       �v:_Fr*@W             c@                           @$3sp@S           P�@������������������������       �e��q.a@E            �[@������������������������       �~��Y@           �{@                            �?	\m1{@�           ��@                          �7@%l#�GX@           �z@������������������������       ���%&�l@�            �j@������������������������       �;)�6��@�            @k@                          �9@{Y�)!@�             w@������������������������       �z�[�d�@�             p@������������������������       �����/@G            �[@�t�b��
     h�h5h8K ��h:��R�(KKKK��h��B�        5@     `r@     Ё@      <@     �I@     �|@     �Z@     �@     `j@     p�@     �v@      C@      2@     �k@     @v@      1@      A@     �s@     �S@      v@     �d@     �v@     �m@      ?@      �?      Q@     �W@              @     �U@      @     `b@      ?@     �a@     �K@      @      �?      I@      T@              @     �Q@      @     �U@      9@     @X@     �F@      @              <@     �J@              @     �G@      �?     �S@      4@     �R@      @@      @      �?      6@      ;@               @      7@       @      @      @      7@      *@                      2@      ,@               @      1@      �?     �N@      @     �F@      $@                      @       @               @      �?              2@              3@      �?                      .@      @                      0@      �?     �E@      @      :@      "@              1@     @c@     `p@      1@      ;@      m@     �R@     �i@     �`@      l@     �f@      <@      *@      a@     �l@      1@      ;@     @h@     @P@     @g@     �\@     �j@     @d@      .@              7@      M@      @      @      N@      @      O@     �@@     �J@     �J@      @      *@     �\@     �e@      ,@      4@     �`@      M@      _@     @T@     �c@     @[@      (@      @      1@      @@                      C@      $@      5@      4@      *@      5@      *@              @      1@                      @      @      �?      $@       @      @      @      @      &@      .@                      ?@      @      4@      $@      @      0@      "@      @      R@     �j@      &@      1@     `a@      ;@     ؃@      G@     �y@     �_@      @             �@@      \@      @      "@     �K@      @     �z@      ,@      j@      G@       @              @      H@              @      4@             �g@      �?     @S@      1@       @              @      0@                       @              `@              F@      @                              @@              @      (@             �M@      �?     �@@      $@       @              =@      P@      @      @     �A@      @     �m@      *@     �`@      =@                      "@      8@                      @      @      A@      @      9@      @                      4@      D@      @      @      =@      �?     `i@      $@     �Z@      7@              @     �C@     �Y@      @       @      U@      6@     @j@      @@     �i@     @T@      @              <@     �O@      @      @      A@      .@     �Z@      6@     �[@     �F@                      0@     �A@      @              0@      "@     �R@       @      C@      ,@                      (@      <@              @      2@      @      @@      ,@     @R@      ?@              @      &@     �C@      @      @      I@      @      Z@      $@     �W@      B@      @      @       @      A@      �?              ?@      @     @R@      @     �O@      ?@      @              @      @      @      @      3@      �?      ?@      @      @@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @i�C%"@�	           ��@       	                     �?��˥��@f           �@                          �5@�/�%�@�            �@                           �?�7�m��@�            �q@������������������������       ���Q��@:            @U@������������������������       ��x/<�@x            �h@                           �?��C�h�	@�            �v@������������������������       ��~~�@=            �\@������������������������       �}�c�ݻ	@�             o@
                           �?���S�@�           ��@                           �?�����@}           ��@������������������������       �lo!�i�@�             k@������������������������       ���y�C^	@�            `v@                           �?��Mq��@R            �@������������������������       ����P�@�            �l@������������������������       ��e?��T	@�           ؆@                            @p�	�_�@L           �@                          �6@���z7�@�           �@                           �?���@fl@�           |�@������������������������       �����N&�?           �x@������������������������       �*�a���@�           ��@                           �?����@
           �y@������������������������       ��ܩ�i@z            �g@������������������������       ��h�@�            �k@                           @�'�ɕ�@�            �p@                           @����I�?f             d@������������������������       ��ט�)� @.            �S@������������������������       ��oc���?8            �T@                           �?kuA@B            �Z@������������������������       �-���L@"             L@������������������������       �����@             �I@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      t@      �@      8@      K@     �z@      T@     Ȑ@      m@     h�@     �t@      >@      .@     �k@     t@      2@      F@     �r@     �O@     0y@     �h@     �u@     `l@      <@      @      L@     �W@      �?      ,@     @V@      5@     @^@     �M@     @[@     �N@      0@              ,@      H@              �?     �C@      @     �P@      3@     �L@      <@      @              @      $@              �?      @      �?      8@       @      <@      (@                      &@      C@                     �A@      @      E@      1@      =@      0@      @      @      E@      G@      �?      *@      I@      .@     �K@      D@      J@     �@@      (@              @      "@              @      *@      @      9@      &@      <@      @      @      @      B@     �B@      �?      @     �B@      (@      >@      =@      8@      :@      @      (@     �d@     `l@      1@      >@      j@      E@     �q@      a@     �m@     �d@      (@      @     �L@     �U@      @      ,@     �T@      *@     �Y@     �H@     �T@     �Q@       @              6@      9@      �?      @     �A@              K@      2@     �C@      0@              @     �A@      O@      @       @      H@      *@      H@      ?@      F@     �K@       @      @     �Z@     �a@      &@      0@     �_@      =@     �f@      V@      c@     �W@      $@              ;@      8@              �?      =@      �?     �P@      *@      G@      5@      �?      @      T@      ]@      &@      .@     @X@      <@     �\@     �R@     �Z@     �R@      "@       @      Y@     �k@      @      $@     �_@      1@     ��@      B@     @{@     @Z@       @       @     �V@     �h@       @      @      ]@      ,@     ��@      ?@      v@     �U@       @              I@      `@       @      @     �S@      "@     �|@      $@     �n@     �O@      �?              $@     �M@              �?      2@             @j@       @      U@       @                      D@     �Q@       @      @      N@      "@     `o@       @     @d@     �K@      �?       @      D@     @Q@              �?      C@      @      Z@      5@      [@      7@      �?       @      >@      <@              �?      .@      �?     �E@      @     �J@      "@      �?              $@     �D@                      7@      @     �N@      .@     �K@      ,@                      $@      9@      @      @      &@      @     �Z@      @     �T@      3@                      @      *@                       @      @     @R@      @      L@       @                      �?      (@                      @      @     �@@              6@      �?                       @      �?                       @              D@      @      A@      �?                      @      (@      @      @      @             �@@       @      :@      1@                      @      @       @       @                      4@       @      *@      @                      @      @       @      �?      @              *@              *@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ"�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���t�@�	           ��@       	                   �5@C�r��@v           Р@                           �?��o^ȣ@�           �@                           �?+E���K@�            �t@������������������������       �k��;�@l             e@������������������������       ��pi��Q@o            �d@                           @r��Af?@�           ��@������������������������       �2�*ֽ@/           �}@������������������������       ���0{��@�             k@
                           �?���5w1	@�           ��@                           �?kv���`	@<           Њ@������������������������       �^��tT@�             l@������������������������       ����R�	@�           ȃ@                           @?�@�            �p@������������������������       �C����@i             e@������������������������       ���81��@=             Y@                           @0�����@L           ��@                           @ڰ�B@<           $�@                           @�"s0�i@�           �@������������������������       �
�����@�           ��@������������������������       ���~�m�@*           P~@                          �5@��;�@B           ��@������������������������       ��/��@�            �r@������������������������       �۽�R�>@�            �l@                           @���zN@             8@������������������������       ��7���� @             &@������������������������       ����G @	             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B 
        4@     r@     �@      6@      H@     p~@     �T@     �@     �g@     p�@     �v@      9@      2@     `j@      s@      0@     �E@     �t@     @P@     �v@     `c@     �w@     �n@      7@      @     �R@     �_@      @      2@     `b@      :@     �o@     @P@     �h@     �X@      @              ?@     �D@      �?      @      <@      @     @\@      .@      S@      0@      @              *@      2@      �?      @      .@      @     @P@      *@      9@       @      @              2@      7@              �?      *@              H@       @     �I@       @              @      F@     @U@      @      ,@     �]@      6@     �a@      I@     �^@     �T@      @      @      5@      K@      @      $@     �S@      1@     @X@      B@     �W@     �N@              @      7@      ?@      �?      @      D@      @     �E@      ,@      ;@      5@      @      (@      a@     @f@      $@      9@     �f@     �C@      \@     �V@     �f@     �b@      0@      (@     @Z@     �`@      $@      2@     �b@     �@@     �P@     �R@     �^@     �]@      ,@      �?      @@      D@      �?      @      D@              =@      "@      C@      <@      @      &@     @R@     @W@      "@      ,@     �[@     �@@     �B@     �P@     @U@     �V@      &@              ?@     �F@              @      ?@      @      G@      .@     �L@      =@       @              @      5@              @      6@      @      C@       @      E@      4@      �?              8@      8@              �?      "@       @       @      @      .@      "@      �?       @     �S@     @n@      @      @     �c@      1@     Є@     �@@     @{@     �\@       @       @     �Q@     @n@      @      @     �c@      (@     Ȅ@      >@      {@     @\@       @       @     �G@     `e@              @     �Y@      @     �@      .@     @r@      P@       @       @      4@     �W@              @     �P@      @     �t@      &@     �d@      :@                      ;@     @S@                      B@             �e@      @     �_@      C@       @              7@     �Q@      @       @      K@      @      d@      .@     �a@     �H@                      $@     �F@      @       @      3@             �^@      @     �S@      ,@                      *@      :@      @             �A@      @     �C@      (@     �O@     �A@                       @                              @      @      �?      @       @       @                      �?                               @      @              @      �?                              @                              �?      �?      �?              �?       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@C��{��@�	           ��@       	                    @���@O           L�@                           �?������@�           $�@                            �?��Ow�@�            �x@������������������������       �𐝾��@F            �^@������������������������       �n��a:�@�            �p@                          �2@�q/�!�@�           �@������������������������       �5V8�i@�            �q@������������������������       �\*��h	@           �z@
                           �?�X��#@�           t�@                            �?�^��Ui @�            �x@������������������������       �Q�)S:��?5            @V@������������������������       �-	��D@�            0s@                          �4@v,	�L@�           ��@������������������������       �3١���@k           ��@������������������������       ��L@J            �^@                           �?��M���@D           ��@                          �7@����@�           ��@                           @���n2�@�            `p@������������������������       �@�k@U            @a@������������������������       �d��៸@M             _@                           @q9~#�@4           �~@������������������������       �(`�p@�             w@������������������������       �"WDTQ@I            @_@                           @7elO		@n           p�@                           �?�HT�E�	@�           H�@������������������������       �:4V�L�@c            `b@������������������������       �AS��r�	@G           `@                          �:@� ����@�            Pr@������������������������       ��P���i@�            �i@������������������������       �i��]?�@;            @V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     h�@     �@@      R@     �z@     @T@     p�@     `j@     x�@     �x@     �A@      @      `@     �s@      "@     �A@      j@      ;@     x�@     �X@     �~@     �g@      0@      @     �T@     @c@      @      8@     �b@      .@      m@     @S@     `k@     �]@      &@              @@     �M@              @      ?@             �Z@      2@     �Z@     �@@      �?              @      8@              �?       @              C@      �?     �D@      @                      <@     �A@              @      7@             @Q@      1@     �P@      <@      �?      @     �I@     �W@      @      4@     @]@      .@     �_@     �M@      \@     �U@      $@      �?      9@     �H@      �?      @      E@      @     @P@      9@      C@      9@      �?      @      :@      G@      @      0@     �R@      &@     �N@      A@     �R@     �N@      "@             �F@     @d@       @      &@     �N@      (@     `|@      5@     q@     �Q@      @              ,@     �K@               @      1@       @     `i@       @     �T@      3@                               @                      �?             �M@              ,@      @                      ,@     �G@               @      0@       @      b@       @      Q@      (@                      ?@     �Z@       @      "@      F@      $@     `o@      3@     �g@      J@      @              =@     @V@       @      "@      ?@      @      l@      2@     �a@     �G@                       @      2@                      *@      @      :@      �?     �H@      @      @      ,@      e@      n@      8@     �B@      k@      K@     �s@     @\@     0r@     `i@      3@       @     �P@      [@      "@      .@     �X@      8@     �a@      C@     �`@     �Z@      "@              =@     �I@      @      @     �D@      @     �M@      @     �A@      6@      @              2@      >@       @       @      9@      @      1@      @      *@      0@      @              &@      5@       @      �?      0@      @      E@              6@      @               @     �B@     �L@      @      (@      M@      2@     �T@      @@     �X@      U@      @      @      ;@      G@      @      (@     �D@      *@     �O@      &@     �S@     �P@      @      �?      $@      &@       @              1@      @      4@      5@      4@      2@              @     �Y@     �`@      .@      6@     @]@      >@      f@     �R@     �c@     @X@      $@      @     @U@     �X@      "@      3@     @U@      5@     �W@     �L@     �V@     @R@      $@              3@      7@                      .@              C@      @      >@      &@      @      @     �P@      S@      "@      3@     �Q@      5@     �L@     �I@      N@      O@      @              1@      A@      @      @      @@      "@     �T@      2@      Q@      8@                      @      :@      @              3@      @      Q@      *@      G@      ,@                      &@       @      �?      @      *@       @      ,@      @      6@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJE��3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@|n�6@�	           ��@       	                    �?T�8Zu@�           �@                           �?�L����@d           ��@                           @��{Gf9@�            �n@������������������������       ���A�M@I             X@������������������������       ���)�3��?j            �b@                            @����ݏ@�            r@������������������������       �������@z            �h@������������������������       �My�Y@ @7            �V@
                           �?�HȈ֪@H           x�@                          �2@��6�|@�            s@������������������������       ���Ʈ�[@�            �j@������������������������       �'� ��@A            �V@                           �?M���d�@�           ��@������������������������       �ֻ�p@�            0r@������������������������       �G����@�            �u@                          �;@��^@
           �@                           @���
!�@�           l�@                            �?<"z�	@            ��@������������������������       ��i�x��@�            �v@������������������������       ��P�K��@           �@                          �8@8&��@�           ��@������������������������       ���"�h2@�           �@������������������������       �ʇ��/3@i            �f@                           @�[/1K	@           �z@                           @_�M�	@�            �t@������������������������       �P��*	@�            �m@������������������������       ��&�?J�@<            �X@                            �?h�`�j�@>            @V@������������������������       ��EL�I@"             H@������������������������       ���S�@            �D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     0t@     0�@      7@      K@     @}@     @S@     �@      g@     Ȉ@     v@     �D@      @      R@     �g@      �?      @     �`@      (@     �@     �O@      w@      [@      @              5@     �M@               @     �@@      @     �m@      &@     �a@      9@                      @     �@@                      2@      @     �]@      @      K@       @                       @      2@                      &@      @     �@@      @      2@      @                      @      .@                      @             @U@              B@      @                      .@      :@               @      .@             @^@      @      V@      1@                      &@      5@                      $@             �T@      @      L@      *@                      @      @               @      @             �C@              @@      @              @     �I@     @`@      �?      @     �Y@      "@     0q@      J@     @l@     �T@      @      @      B@      A@      �?       @     �F@      @      D@      A@     �K@      F@      @      @     �@@      :@                     �C@       @      7@      8@     �C@      8@      �?       @      @       @      �?       @      @      @      1@      $@      0@      4@      @              .@      X@              @     �L@      @     `m@      2@     `e@     �C@                      @      F@                      B@             �\@      $@     @P@      1@                      $@      J@              @      5@      @     @^@       @     �Z@      6@              ,@     `o@     �v@      6@     �G@     �t@     @P@     �@     @^@     �z@     �n@     �B@      @      i@     `r@      1@      A@     pp@     �I@      }@      Y@      x@     �d@      >@      @     @d@      g@      *@      <@     @f@      C@     �f@     �S@     `h@     @Y@      <@             �N@     �B@      �?      0@      H@      (@     �L@      ;@     @P@      =@      @      @     @Y@     �b@      (@      (@     @`@      :@     @_@     �I@     @`@      R@      5@      �?     �C@     @[@      @      @     @U@      *@     �q@      6@     �g@      P@       @      �?      @@     �W@      @      @      R@      $@     �l@      @     �a@      E@       @              @      ,@      �?      �?      *@      @      K@      2@      H@      6@               @      I@     �P@      @      *@     �Q@      ,@      H@      5@     �D@      T@      @       @     �E@      H@      @      *@     �I@      *@      ?@      5@      :@     @Q@      @      @      ?@      G@      @      @      B@       @      .@      &@      1@     �H@      @      @      (@       @              @      .@      @      0@      $@      "@      4@                      @      3@                      3@      �?      1@              .@      &@                      @      .@                      �?      �?      $@              "@       @                      @      @                      2@              @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJۛ:-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�&�1k@�	           ��@       	                    �?��O�v�@i           �@                          �<@s[9���@�           �@                          �6@�{�>@z           Ђ@������������������������       �r ϓ@           �z@������������������������       �����@u            @f@                           �?������@,            @R@������������������������       �D� �c@             :@������������������������       ��E��$@            �G@
                           �?Iv���	@�           ��@                           �?�ㆢM
@�           p�@������������������������       ��A]쬆@
           py@������������������������       �;�
�P{
@�           (�@                            @t�!'0Z@           �x@������������������������       ����<@�            �q@������������������������       �w*L��@L            @\@                           @�](�B@7           �@                           @�r��@�           ̒@                           @ڔA��@.           P�@������������������������       �P�JL��@�           ��@������������������������       ��ϔ�
�?L            �]@                          �4@�n�:� @�            �t@������������������������       ����"1�?u            @h@������������������������       �%-iݧI@S            �`@                            �?����@A           @�@                          �5@�ĥ�;�@M            ``@������������������������       ����^� @,            �Q@������������������������       ��d�T@!            �N@                           �?�0�>��@�            Px@������������������������       ��b+��v@Z            �a@������������������������       ���&U!*@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     0p@      �@      ;@     �P@     �|@     �V@     ��@      n@     ��@     �w@      =@      4@     @h@     �t@      4@     �I@     �s@     �M@     �w@     �h@      u@     �o@      :@      �?     �Q@     @W@      �?      (@      T@      @      d@     �C@     �b@      P@      @      �?      N@     �T@      �?      "@     �Q@      @     �c@      ?@      a@      G@      @              D@      L@              @      B@      �?      ^@      ;@     �Y@     �A@      �?      �?      4@      :@      �?      @     �A@       @     �C@      @      A@      &@       @              &@      &@              @      "@              �?       @      (@      2@                      "@      @                      @              �?              @      @                       @       @              @      @                       @      "@      &@              3@     �^@     �m@      3@     �C@     �m@      L@     �k@      d@     �g@     �g@      7@      3@      Y@     �d@      1@      @@     �d@     �G@     @b@      ^@     �_@      c@      7@      �?      4@     �R@      @      1@     �P@       @     �P@     �A@     �I@      M@      @      2@      T@      W@      *@      .@      Y@     �C@     �S@     @U@      S@     �W@      2@              7@     �Q@       @      @     @Q@      "@      S@      D@     �O@     �C@                      2@     �E@              @     �M@      @     �H@      ;@     �J@      9@                      @      <@       @              $@      @      ;@      *@      $@      ,@                     @P@     �j@      @      .@     @b@      @@     ��@     �D@     @|@     @^@      @              D@     �c@       @      @     �Y@      ,@     �}@      4@     @s@     �S@       @              A@      X@       @       @     @V@      ,@     �t@      2@      l@      O@       @              ?@      W@       @       @     @R@      ,@     @q@      2@     �g@      L@       @              @      @                      0@             �K@              A@      @                      @      N@               @      ,@              b@       @      U@      0@                       @      ;@               @      @             �Y@              H@      @                      @     �@@                      @              E@       @      B@      &@                      9@      M@      @      &@     �E@      2@     �b@      5@      b@     �E@      �?              @      @      �?      �?      .@       @      G@      @     �@@      @                      �?       @              �?      &@             �A@      �?      ,@      @                      @      @      �?              @       @      &@      @      3@       @                      2@     �I@      @      $@      <@      $@     @Z@      .@     �[@      B@      �?              @      3@              @      @              K@      @      E@      @                      &@      @@      @      @      8@      $@     �I@      &@     @Q@      =@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��a��I@�	           ��@       	                    �?lhվ��@v           \�@                           �?�@P!	@
           ��@                          �5@���}��@7           �}@������������������������       ��B�9@�             n@������������������������       �ui���@�            �m@                          �5@_�~?��	@�           (�@������������������������       �ĕ�k�%@G           ��@������������������������       ��UV�R
@�           ��@
                           �?[��-@l           0�@                            �?���@s             g@������������������������       �^6rF%@&            �P@������������������������       �N웇Â@M            �]@                           �?-hҊ��@�            �x@������������������������       �UO!@             :@������������������������       �v{W��q@�            0w@                          �7@�}�j�@3           l�@                           @:c���@/           ��@                           �?P~0���@�            �s@������������������������       ��ue!�?@c            @d@������������������������       �<L�" @`             c@                          �4@>
�P�@l           �@������������������������       ��6�@�           �@������������������������       �m0��~�@�            r@                            �?%z��>@           �y@                           @Q:�� @�             j@������������������������       �ɱ%(�@;            �S@������������������������       �X`�jQ@P             `@                           �?h��A��@y            �i@������������������������       ����1�@6            �V@������������������������       ��͖~t�@C             ]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     �r@     H�@      A@      G@      ~@     �U@     ��@     �k@     h�@     0v@     �@@      &@     @m@     �t@      8@      C@     �t@     @P@     @y@      g@     �t@     �m@      <@      &@     �f@     `o@      8@      <@     Pp@     �G@      o@      b@     `m@     �f@      9@              J@     @T@              $@      R@      @     �W@      5@      Y@      E@      �?              .@     �B@              @      >@      @     @S@       @      J@      ,@      �?             �B@      F@              @      E@      �?      2@      *@      H@      <@              &@     ``@     @e@      8@      2@     �g@     �E@      c@     �^@     �`@     �a@      8@      @     �I@      W@      @      @     �U@      $@     @Y@     �H@     �R@     �J@      @       @      T@     �S@      4@      ,@     �Y@     �@@      J@     �R@      N@      V@      1@             �I@      T@              $@     �Q@      2@     �c@     �D@     �X@     �K@      @              (@      0@              �?      6@       @      R@      @      F@       @       @               @      "@              �?      @              5@              8@      �?       @              $@      @                      .@       @     �I@      @      4@      @                     �C@      P@              "@      H@      0@      U@     �A@      K@     �G@      �?               @      �?              @       @      �?      �?      $@              @                     �B@     �O@              @      G@      .@     �T@      9@      K@     �E@      �?             @Q@     �k@      $@       @     �b@      5@     ��@      B@      |@     @]@      @             �F@     �e@      @       @     @V@      ,@     �@      3@      u@     �R@      @              1@     �J@                      .@      &@     �^@       @     �P@      2@      @              *@      5@                      &@      @      H@      @      B@      .@      @              @      @@                      @      @     �R@      �?      ?@      @                      <@     @^@      @       @     �R@      @     px@      &@     �p@      L@      �?              ,@      S@      @       @      E@             �r@      @     @h@      B@      �?              ,@     �F@       @              @@      @     �W@      @     �R@      4@                      8@      H@      @      @      O@      @     �V@      1@      \@     �E@                      .@      =@              �?      3@      @     �G@      *@     �L@      5@                       @      &@                      @      @      0@      @      3@      *@                      *@      2@              �?      (@       @      ?@      @      C@       @                      "@      3@      @      @     �E@      �?      F@      @     �K@      6@                      @      ,@               @      2@              6@      �?      5@      @                      @      @      @      @      9@      �?      6@      @      A@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��uhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��LT,`@�	           ��@       	                    �?VI��b@�           ��@                           �?g���@$           p}@                            @ ^40@h            �e@������������������������       ���}�ب@F            @^@������������������������       ��j���m@"             J@                            �?�j?ׁ�@�            �r@������������������������       � �2��!@Y            @b@������������������������       �О�z�@c             c@
                           @�++�b�@�           @�@                          �2@���� @]           h�@������������������������       ��#�5P�?�            �m@������������������������       ��Si@.@�             t@                            @<�>4�@v            `g@������������������������       �c�7ȓ�@_            @c@������������������������       �=*,I�R @            �@@                          �6@�'?D@�           �@                           @�; ӓ4@           0�@                          �1@�$qMN�@�           ܐ@������������������������       �����ۥ@�            �o@������������������������       �'=�AG@           ؉@                           @?���@\           ��@������������������������       �M�Փ@�            u@������������������������       ��o"1X�@�            �h@                            @���W�>	@�           ��@                           @(�R���@�           ��@������������������������       ����)�z	@           py@������������������������       ����E�@�            �s@                           @5����	@�            �v@������������������������       �=d&n�
@�            �q@������������������������       ��M�VM6@1            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@      t@     ��@      =@     �L@     �|@     @W@     �@     �i@     0�@     �u@      ?@             �R@     �f@      @      0@      W@       @     p{@     �B@     �q@     @S@      @             �F@     @U@       @      $@      K@       @     �V@      :@     @Z@     �G@      @              5@      ?@                      0@             �D@       @     �H@      (@      �?              .@      3@                      ,@              9@      �?      A@      (@      �?              @      (@                       @              0@      �?      .@                              8@      K@       @      $@      C@       @      I@      8@      L@     �A@      @              $@      7@      �?      @      .@              2@      1@      ;@      9@      @              ,@      ?@      �?      @      7@       @      @@      @      =@      $@                      >@     �W@       @      @      C@      @     �u@      &@     @f@      >@                      6@      R@              @      ;@      @     0q@       @     �`@      2@                      @      ?@                      &@             �a@             �F@      @                      2@     �D@              @      0@      @     �`@       @     �U@      *@                       @      7@       @       @      &@      �?     @R@      "@      G@      (@                      @      7@       @              @      �?      M@      "@     �B@      $@                      �?                       @      @              .@              "@       @              .@     �n@     �w@      9@     �D@     �v@     @U@     0�@      e@     X�@     �p@      ;@      @     �_@     @l@      0@      8@      k@      B@      x@      T@     @v@     �`@      @      @      U@     �`@      *@      0@     @c@      6@     `p@      E@     �p@     @U@                      0@      ;@              �?      6@             @T@      (@      S@      1@              @      Q@     �Z@      *@      .@     �`@      6@     �f@      >@     �g@      Q@               @      E@     @W@      @       @      O@      ,@      _@      C@      W@     �H@      @       @     �A@     �Q@       @      @      I@      (@      K@     �B@     �C@      9@      @              @      6@      �?      @      (@       @     �Q@      �?     �J@      8@      �?      "@     @^@     `c@      "@      1@     �b@     �H@     �`@      V@     �h@      a@      5@      @     @R@     �W@      @      "@      X@      @@     �S@      Q@     �b@      Y@      *@       @      G@     �F@      @      @     �M@      8@      ;@      K@     �P@      N@      *@      �?      ;@      I@              @     �B@       @      J@      ,@     �T@      D@              @      H@      N@      @       @      K@      1@     �J@      4@     �H@      B@       @      @     �F@     �J@      @      @      C@      0@      @@      3@      ;@      =@       @              @      @              �?      0@      �?      5@      �?      6@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ13�jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��}��@�	           ��@       	                    �?�(M�D	@h           <�@                          �8@���@�@�           ��@                          �5@�ͧ�@%           �~@������������������������       �4DM��@�            pv@������������������������       �[��*@N            �`@                          �?@A���/@e            �d@������������������������       �`)��@X             b@������������������������       ���[^D@             4@
                           �?(İ%��	@�           8�@                           �?��J�s+
@�           ��@������������������������       �`� ́
@�            �x@������������������������       ��E-��	@�           ��@                          �4@|�P�+@           �z@������������������������       �� �"%@�             g@������������������������       �`%0
�@�            @n@                            �?�و\͕@8           ��@                           @Vؖ��<@�             x@                          �3@g%Q5��@@            @[@������������������������       ��:0���?              N@������������������������       �)%�Ha\@             �H@                          �6@��6d-�@�            0q@������������������������       �c.���h�?}            `h@������������������������       �Z���~@5             T@                           @�� b�@F           ��@                            @sK?���@I           H�@������������������������       ��&�B@�           ��@������������������������       �� [K�?�?`            �b@                           �?�M"H,�@�             x@������������������������       �_�"��@_            �`@������������������������       �G���At@�            �o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     s@      �@      A@     �O@     �z@     �T@     ��@     �l@     ��@     `v@      C@      6@     �m@     �u@      9@      J@     Pr@     @P@     0v@     @h@     u@     @n@     �@@       @     �P@     @]@      �?      (@     �Q@      @      c@      =@     ``@     �N@      @              K@     @T@      �?      @      F@      @      `@      7@     �[@      C@       @              =@     @P@      �?      @      7@      @     �X@      3@      U@      :@       @              9@      0@                      5@              =@      @      :@      (@               @      *@      B@              @      ;@      @      8@      @      5@      7@      @       @      @     �@@               @      6@      @      8@      @      5@      6@      @              @      @              @      @                      �?              �?              4@     @e@     @m@      8@      D@     �k@      M@     `i@     �d@     �i@     �f@      ;@      4@     @`@     �e@      4@      ?@      e@     �F@      ]@     �_@     �`@     ``@      :@       @      F@     @R@      $@       @      J@      2@      L@      D@      <@      I@      $@      (@     �U@     @Y@      $@      7@     @]@      ;@      N@     �U@     �Z@     @T@      0@              D@      N@      @      "@     �J@      *@     �U@     �C@     �Q@      I@      �?               @      :@      @              :@       @     �K@      3@      <@      1@                      @@      A@              "@      ;@      &@      @@      4@     �E@     �@@      �?              Q@     �l@      "@      &@     �`@      1@     x�@     �A@     �z@      ]@      @              &@     �E@      �?      �?      3@      @     �f@      .@     �R@      @@                      @      3@                      �?              I@      @      (@      .@                              @                                     �A@      @      @      "@                      @      ,@                      �?              .@       @      @      @                      @      8@      �?      �?      2@      @     �`@       @     �O@      1@                      �?      @              �?      (@       @     �]@      �?      F@       @                      @      1@      �?              @       @      ,@      @      3@      "@                     �L@     @g@       @      $@     �\@      *@     �}@      4@      v@      U@      @              E@      `@       @      @     �S@      @     Pw@      @     �m@     �I@      @             �A@     �^@       @      @     �P@      @     �r@      @      h@     �H@       @              @      @                      (@             �R@      �?     �G@       @      �?              .@      M@      @      @     �A@      @     �X@      *@     �\@     �@@       @              @      1@                       @             �J@      @      D@      @       @              (@     �D@      @      @      ;@      @      G@       @     �R@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJtz+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@>���Y@�	           ��@       	                    @TG2rDC@           Ȝ@                           �?{�)S@7           0�@                           �?;8vN�@�           ��@������������������������       ��~ �}�@y            �h@������������������������       �2\�s@	           �z@                            �?�V�Y�@�            `q@������������������������       �#�nFy@6            �U@������������������������       �o"+0�@            �g@
                           @�\,;@H           `�@                          �1@�Ӈ�8@�            �l@������������������������       �� ;ɳM @>            �[@������������������������       ��!���@J            �]@                           �?�6��@�           8�@������������������������       ����D�@�            v@������������������������       ��^k!<@�            `v@                            �?/{� a�@           .�@                           @��W�@�           8�@                          �<@�!��J@f           ��@������������������������       ��h�k��@           Љ@������������������������       ��J��@b            �c@                          �5@;��%�h@J             ^@������������������������       ��D����@
             *@������������������������       ��S�Z1X@@            �Z@                           �?���d@i           H�@                           �?S��*�	@(           �}@������������������������       �`z��@C            @Z@������������������������       �Ùm��	@�            w@                           @�?$��@A           �~@������������������������       ��q��Z�@           �{@������������������������       ��	�@$            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     `s@     ��@      A@      L@     P|@      R@     ��@     �m@     ��@     �u@      ;@      @      ]@     `o@      @      ,@      e@      &@      �@     �Z@     �w@     @`@       @      @     @Q@      a@      @      "@     �[@       @      m@     �U@      b@     �U@      @      @      I@     @V@       @       @     �U@       @     �a@      O@     �W@     �Q@      @              $@      A@               @      (@       @     �L@      .@      C@      <@      �?      @      D@     �K@       @      @     �R@      @     @U@     �G@      L@      E@      @              3@      H@      @      �?      8@             �V@      9@      I@      1@                      @      ,@                      @              <@       @      <@      @                      .@      A@      @      �?      2@             �O@      7@      6@      (@                     �G@     �\@       @      @     �M@      @     py@      4@     �m@     �E@      �?              5@     �C@                      "@      @     @U@      @     �J@      ,@                      @      &@                      @             �J@      �?      =@      @                      ,@      <@                      @      @      @@      @      8@      "@                      :@     �R@       @      @      I@              t@      .@     @g@      =@      �?              @      ?@       @      @      :@             �c@       @      X@      3@                      3@      F@                      8@             `d@      @     �V@      $@      �?      .@     @h@     Ps@      ;@      E@     �q@     �N@      w@      `@     `y@      k@      3@      @     @_@     �b@      *@      9@      a@     �@@     �h@     �T@      l@      Y@      "@      @      Z@     �`@      (@      8@     @_@      8@     @g@     �K@     �j@     �W@       @      @     �V@      ]@      (@      4@     �[@      .@     �e@      B@     �g@     �I@      @              *@      0@              @      ,@      "@      &@      3@      8@      F@       @       @      5@      1@      �?      �?      &@      "@      &@      <@      *@      @      �?      �?              @              �?      �?      @      �?                      �?              �?      5@      *@      �?              $@      @      $@      <@      *@      @      �?       @     @Q@      d@      ,@      1@     �b@      <@     `e@      G@     �f@     @]@      $@      @     �C@     �W@      &@      .@      S@      4@     �E@      ?@     �P@     @P@      @              @      <@      @      @      0@              .@       @      4@      @              @      A@     �P@       @      (@      N@      4@      <@      7@      G@      M@      @      �?      >@     �P@      @       @      R@       @      `@      .@     �\@      J@      @      �?      8@      J@      @       @      N@      @     �^@      *@     @Z@      J@                      @      ,@                      (@       @      @       @      $@              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�%��
}@�	           ��@       	                    �?���k�5@           D�@                            @��u@F�@.           ~@                           �?=�ߓ�@�            �q@������������������������       ��ݪp�c@S             `@������������������������       ����W�@b             c@                           �?�f0���@y            �h@������������������������       �e
��?$            �P@������������������������       ���$R�=@U            �`@
                          �5@��1?�@�           ��@                            �?7Գ�!*�?N           x�@������������������������       �C壋�E @�            �q@������������������������       �!G\v�h�?�            �n@                          �8@(A�w�@�             l@������������������������       �\��]g8@M            �\@������������������������       ���o#G@D            �[@                           @�bc��t@�           �@                           �?����	@�           �@                          �<@���Y�	@�           ��@������������������������       ���+��	@\           ��@������������������������       �8,�'	@_            �b@                           �?�V����@           0y@������������������������       ��+�㣅@             B@������������������������       �a7:�fq@�            �v@                           @k�J�?�@�           �@                           @���I@�           ��@������������������������       ��*��b�@�            �n@������������������������       ��[�	��@U           �@                          �3@�S�yE�@�            @v@������������������������       �萧%P@F             \@������������������������       �~�y�@�            �n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      @@      N@     0~@      X@     H�@     @k@     (�@     @u@      @@             �Y@     `e@      �?      (@     @W@       @     �|@      @@     �p@     �S@      @             �Q@     �T@              "@      K@      @     �Z@      2@     @V@     �G@      @             �G@     �D@               @      B@       @      J@      $@      L@     �@@      @              3@      *@                      0@              A@      @      ;@      .@       @              <@      <@               @      4@       @      2@      @      =@      2@      �?              7@     �D@              @      2@      �?      K@       @     �@@      ,@                      @      *@                      @              <@              2@                              3@      <@              @      ,@      �?      :@       @      .@      ,@                     �@@     @V@      �?      @     �C@      @     @v@      ,@     `f@      ?@       @              0@     �O@              @      9@      �?     �q@      @      ^@      $@                      "@     �F@              @      .@      �?      b@      �?      L@       @                      @      2@                      $@              a@      @      P@       @                      1@      :@      �?              ,@      @     �R@      @     �M@      5@       @              .@      *@      �?              "@              C@       @      9@      &@                       @      *@                      @      @      B@      @      A@      $@       @      4@      h@     px@      ?@      H@     `x@      V@     ؀@     @g@     �@     `p@      ;@      3@     �`@     �m@      5@      ?@     pp@      Q@      i@     �c@     @j@      e@      7@      3@      [@      d@      4@      6@     `i@     �L@     �`@     �Y@     @b@      a@      6@      2@     �U@     �a@      0@      4@     �f@      F@     �_@     @V@     @`@     �Z@      5@      �?      5@      3@      @       @      7@      *@      @      ,@      0@      =@      �?              9@      S@      �?      "@      N@      &@     @Q@     �K@      P@      @@      �?              @      "@              @      @              �?      @      @      @                      6@     �P@      �?      @      K@      &@      Q@      I@     �N@      ;@      �?      �?      N@     @c@      $@      1@     �_@      4@      u@      <@     pr@     �W@      @      �?      B@     �\@       @      @     �S@      @     @p@      3@     @k@      I@       @      �?      1@     �C@       @              4@      @     �R@      @      L@      6@      �?              3@      S@              @      M@              g@      (@     @d@      <@      �?              8@     �C@       @      *@     �H@      *@     �S@      "@     @S@      F@       @              @      (@      �?      @      $@              E@       @      :@       @                      3@      ;@      @      @     �C@      *@      B@      @     �I@      B@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>��MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@q(��x@�	           ��@       	                    �?j�=�@�            �@                          �2@���3j@^           ��@                           @�>�Q�?@           y@������������������������       �쎕72x@w            `d@������������������������       �P1?����?�            �m@                           @*	�� @P            �_@������������������������       ����#l@0            @Q@������������������������       ����|���?              M@
                           �?�^��@(           ��@                           @[�nW@�            s@������������������������       �x����@�             q@������������������������       �y�^���@             ?@                          �1@\_�+�@k           8�@������������������������       �G/���1@�            �n@������������������������       �`���(�@�            u@                           �?"����@           ��@                           �?XS�b@�           H�@                          �<@��=��@�             t@������������������������       ��IHy0@�            pp@������������������������       ��͸ 2�@%            �L@                           �?&��h��@�            �x@������������������������       ����#�J@�            @m@������������������������       ���Pz@k            �c@                           @�%x %	@U           ��@                            @nY��	@3           �@������������������������       ��KwoV�@�           �@������������������������       �qM��;	@[           ��@                           �?0,�r@"            �J@������������������������       �,�\;� @             4@������������������������       �rc��r@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �t@     H�@      <@     �N@     0}@      U@     0�@     �i@     h�@     �u@     �@@      @      R@     �f@      @       @     �[@      *@     �@      L@     u@      _@       @              6@     �J@               @      <@      �?     �l@      *@     `c@      6@      �?              3@      F@               @      8@             �g@       @     @X@      .@      �?              ,@      1@              �?      1@              L@      @     �F@      "@                      @      ;@              �?      @             �`@      @      J@      @      �?              @      "@                      @      �?      D@      @      M@      @                      @      @                      @      �?      ,@      @      >@      @                              @                      �?              :@              <@                      @      I@     �_@      @      @     �T@      (@     q@     �E@     �f@     �Y@      �?      @      ;@      C@       @      @     �F@      @     �H@      >@     �I@      H@      �?      @      7@     �A@       @      @     �B@      @     �G@      <@      F@      H@                      @      @                       @      @       @       @      @              �?              7@     @V@      @      @      C@      @      l@      *@     ``@      K@                      @      D@               @      @             �\@      @     �I@      4@                      0@     �H@      @      �?      ?@      @     @[@      "@      T@      A@              5@      p@     Pw@      7@     �J@     @v@     �Q@     �~@     �b@     �{@      l@      ?@      �?      O@     @[@              .@     �R@      &@      k@      1@      b@     �I@      $@      �?      G@      J@              $@      G@      �?      J@      (@     �J@      C@      "@      �?      D@      F@              @      C@      �?      I@      &@     �I@      ,@      "@              @       @              @       @               @      �?       @      8@                      0@     �L@              @      =@      $@     �d@      @      W@      *@      �?              "@      A@              @      4@      @     �[@       @     �D@      @                      @      7@                      "@      @      K@      @     �I@      @      �?      4@     �h@     �p@      7@      C@     �q@      N@     Pq@     ``@     �r@     �e@      5@      1@     `g@     `p@      4@      C@     �p@      M@     �p@     �^@     �r@     �e@      2@      $@      _@      d@      @      <@     �e@      E@     @i@      U@      j@     �Z@      &@      @     �O@     @Y@      ,@      $@     @W@      0@     @Q@     �C@     �V@     @P@      @      @      "@       @      @              ,@       @      @       @      �?       @      @      @       @      �?                      @              �?      @      �?              @              @      �?      @              $@       @      @      @               @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ7^8RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @I>���u@w	           ��@       	                    �?8M0 	@I           ��@                           �?2r��G	@            �@                           �? ^S)z�@�             s@������������������������       �Sj��k@�             k@������������������������       ��^�=��@7            �V@                            �?��S=��	@J           p�@������������������������       �o�uW_@�            pr@������������������������       �����	@�            pp@
                           �?X���/�@A           Г@                          �7@>��*X�@           �x@������������������������       �̖�&�@�             o@������������������������       ��B�d�@\            `b@                          �4@t�{�	@=           @�@������������������������       �O � @�            �t@������������������������       �P��W�|	@d           ��@                           @�*�^@.           ԛ@                           @S�t��@�           (�@                           @m).���@�            �x@������������������������       ��5��w@�            �r@������������������������       ��xKG!�@;            �X@                            @V�V'�G@�           ��@������������������������       �C�Hqܘ@�           0�@������������������������       �R� ���?9            @V@                          �?@ڄ��Q@O           X�@                            @�dI�@G           Ѐ@������������������������       �	`/sE�@�            0z@������������������������       ���XG�@S            �]@������������������������       ��߆dӚ�?             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �t@     Ђ@     �B@      I@      z@     �W@     (�@     �j@     x�@     �t@     �B@      1@      m@     0u@      @@      ?@     �q@     @S@     �t@      f@     �u@     `l@      =@       @     @R@     �c@      3@       @     @\@      F@      `@     @S@     @]@     �[@      $@              8@      D@      @      @     �A@       @     �R@      8@     �L@     �A@       @              4@      @@      @      @      8@      @      C@      4@     �C@      =@       @              @       @                      &@      @      B@      @      2@      @               @     �H@      ]@      .@      @     �S@      B@     �K@     �J@      N@     �R@       @              8@     �P@       @      @     �J@      5@      :@     �C@      4@      A@      @       @      9@     �H@      *@      �?      9@      .@      =@      ,@      D@     �D@      @      "@      d@     �f@      *@      7@     �e@     �@@     �i@     �X@      m@     @]@      3@      �?     �Q@      D@              "@      I@      @     @P@      @@      V@      >@       @      �?      E@      7@              @      ;@             �G@      *@     �Q@      6@                      <@      1@              @      7@      @      2@      3@      2@       @       @       @     �V@     �a@      *@      ,@     �^@      >@     �a@     �P@      b@     �U@      &@              2@     �E@      @      @      H@      @      U@      3@     @Q@      ?@      @       @      R@      Y@      @      &@     �R@      :@     �L@      H@      S@      L@      @      �?     @X@     pp@      @      3@     @`@      1@     ��@      C@     {@      [@       @      �?     �N@     �e@              @     @T@      $@     �@      .@     0s@     �O@      @      �?      >@      Q@              �?      A@      $@      a@      @     @U@      4@      @      �?      .@      L@              �?      5@      "@     �Z@      �?     @Q@      1@                      .@      (@                      *@      �?      =@      @      0@      @      @              ?@     �Z@              @     �G@              w@      "@     �k@     �E@      �?              >@     @Z@              @     �D@             `t@      "@      g@     �D@      �?              �?      �?                      @              E@             �B@       @                      B@     @V@      @      ,@     �H@      @     �c@      7@     �_@     �F@      @             �A@     @V@      @      ,@     �H@      @     �c@      6@     @_@     �A@      @              A@     @T@      @      "@      E@      �?     @[@      4@     @X@      4@      @              �?       @       @      @      @       @     �H@       @      <@      .@                      �?                                      @              �?      �?      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��Z�@�	           ��@       	                    @��=C�@�           �@                           �?3����@c            �@                          �;@��۰�@           y@������������������������       �WY��m�@�            v@������������������������       ��V�@             H@                          �<@S#I\f	@W           ��@������������������������       �-I�B4	@           8�@������������������������       �Ŝ���@@D             \@
                           @4G�r�F@�           ��@                           @>g(^gf@�           ��@������������������������       �c8	�f@�           \�@������������������������       �̴]E=@             3@                           �?�'��O�@�             x@������������������������       ��~َb�@a            �c@������������������������       ����`<�@�            �l@                           @)���@�           T�@                          �9@�ތ��@"           ��@                           �?��l��@�           P�@������������������������       ��V�3�@�            Px@������������������������       �Ln��R@�            Pr@                          @A@��N@,:@i            `e@������������������������       �8��eH@b            �c@������������������������       ��D=�U�@             (@                          �1@Z��Wg�@�             p@                           �?�j���Q @             ;@������������������������       ��"�@}��?
             .@������������������������       �^�z|�X�?             (@                           @����'	@�            �l@������������������������       ����y�@j            �e@������������������������       �f�r��@!            �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �q@     8�@      8@      F@     �{@     @U@     4�@     �k@     `�@     �v@      :@      *@     `i@     �x@       @      :@     �r@      N@     8�@      d@     p�@      p@      6@      &@     `b@     �g@       @      5@     @h@      H@     �k@      `@     �j@     �b@      0@       @     �I@     �K@              @     �E@      @     �U@      7@     �X@      @@       @             �E@     �I@              @     �D@      @     �U@      0@     @V@      2@       @       @       @      @              �?       @      �?              @      "@      ,@              "@      X@      a@       @      1@     �b@      F@     �`@     �Z@      ]@     �]@      ,@       @     �U@      `@       @      0@      a@      9@      `@     �V@     �[@      W@      $@      �?      $@       @              �?      ,@      3@      @      0@      @      ;@      @       @      L@     @i@              @     �Y@      (@     H�@      @@     �w@     @Z@      @       @     �C@     `a@                     �P@      @      |@      1@     �p@     @R@      @       @      B@     `a@                      P@      @     �{@      &@     �p@     @Q@      @              @                               @      �?      @      @              @                      1@     �O@              @     �B@      @     @Z@      .@     �Z@      @@                       @      9@              @      ,@             �L@      @     �D@      $@                      .@      C@               @      7@      @      H@      $@     �P@      6@              @     �T@     �c@      0@      2@     �b@      9@     `p@     �N@     �k@     �Z@      @      @     �P@     �[@      $@      "@      ^@      .@     �i@      C@     �h@     @S@              @     �H@     �V@      "@      @     �U@      &@     `g@      7@     �d@      J@              @     �C@      J@      "@      @     �P@       @     @P@      3@      V@     �B@                      $@     �C@              @      4@      @     �^@      @     @S@      .@              @      1@      4@      �?      @      A@      @      1@      .@      @@      9@                      ,@      2@              @      @@      @      1@      ,@      @@      9@              @      @       @      �?               @                      �?                                      1@     �G@      @      "@      <@      $@      M@      7@      9@      =@      @              @                               @              ,@      �?       @      @                       @                              �?               @      �?              @                       @                              �?              @               @      �?                      *@     �G@      @      "@      :@      $@      F@      6@      7@      9@      @               @      E@       @       @      4@      "@      ?@      6@      ,@      ,@      @              @      @      @      �?      @      �?      *@              "@      &@        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�Z�<@�	           ��@       	                    �?p�P��6@k           ��@                          �2@G$���@j           ��@                            @k�K�ܪ@�            �u@������������������������       ������@m            �f@������������������������       ��2��?@[             e@                           @e��B��@�            �n@������������������������       �/Ш#�*@|            �h@������������������������       ���C	��@&             I@
                           @��oC@           <�@                           @�糂�.@�            `p@������������������������       ��U�� �@Q             ^@������������������������       ���B2@Z            �a@                            �?��`.2@V           H�@������������������������       �S2��]@L           (�@������������������������       ��?����@
           @|@                           �?��W�d@-           P�@                            �?�N|vR�@�           Ђ@                           �?�}+��\@�            u@������������������������       �[M#ʻY@m            �e@������������������������       �j�}��@g            �d@                           @�@%Y�D@�            �p@������������������������       ��Q�x�2@d             d@������������������������       ���1�F� @H             Z@                          �:@U6W^��@�           8�@                           @$b�u@�           ��@������������������������       ����'	@�           h�@������������������������       �����@�            �x@                           �?tMUkl�@            }@������������������������       �)��~U�@�            �o@������������������������       ������@{            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      r@     @�@      9@      J@      �@     �R@     ��@     `k@     ��@     w@      <@      @     �W@     �l@      &@      $@     �g@      3@     �@     @V@     x@     �a@      &@      @     �E@     �R@       @      @     @[@      (@     @\@      H@     �Z@      Q@      $@      �?      =@     �G@      �?      @     @R@       @     �R@      5@     �O@      @@      �?      �?      4@      :@                      <@             �@@      $@     �F@      0@      �?              "@      5@      �?      @     �F@       @     �D@      &@      2@      0@               @      ,@      <@      �?              B@      $@     �C@      ;@      F@      B@      "@      �?      &@      8@                      =@      $@      >@      1@     �D@      :@      @      �?      @      @      �?              @              "@      $@      @      $@       @             �I@      c@      "@      @     �T@      @     ��@     �D@     `q@     @R@      �?              @      B@      @      @      =@       @     @V@      5@     �J@      3@                      @       @              @      4@      �?     �C@      @      =@       @                      �?      <@      @              "@      �?      I@      .@      8@      &@                      F@     @]@      @      @     �J@      @     �{@      4@      l@      K@      �?              6@      M@      @      @     �A@             `k@      @     �`@     �@@                      6@     �M@                      2@      @     �k@      *@     �V@      5@      �?      0@     @h@     @t@      ,@      E@     t@      L@     0w@     @`@     pw@     �l@      1@             �L@     @Y@       @      "@      R@      @     �b@      =@     �]@      K@      @             �A@     �L@       @      @     �@@      @      Q@      1@      R@     �C@      @              1@      :@      �?      @      3@      @      E@      (@      ;@      5@                      2@      ?@      �?      �?      ,@      �?      :@      @     �F@      2@      @              6@      F@              @     �C@      �?     @T@      (@     �G@      .@                      3@      <@              @     �A@              A@      &@      4@      $@                      @      0@                      @      �?     �G@      �?      ;@      @              0@      a@     �k@      (@     �@@      o@     �I@     �k@     @Y@      p@     �e@      (@      @     �U@      e@      "@      9@      d@      ;@     �d@     @R@     �g@     @X@      (@       @      R@     @]@       @      3@      \@      6@      L@     �L@      T@      Q@       @      �?      .@      J@      �?      @     �H@      @     �[@      0@     �[@      =@      @      *@      I@      K@      @       @      V@      8@      L@      <@     @P@     @S@              *@      5@      6@      @       @     �B@      1@      9@      3@      =@      P@                      =@      @@              @     �I@      @      ?@      "@      B@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ벘=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @.�M�"@�	           ��@       	                   �5@���ᘺ@d           :�@                           @�J�l@�           T�@                           �?��N��o@           ��@������������������������       �����L@i           `�@������������������������       �5�ߑ@�            @r@                          �0@M����	@�            �l@������������������������       �)���	@             1@������������������������       �N�vu�	@�            �j@
                           �?^�W!�|	@�            �@                          �:@	B,�	@
           0�@������������������������       ��h���@	@K           ؀@������������������������       ���]�U	@�            �r@                           �?6b&wt @�             p@������������������������       ��,��@0            @R@������������������������       ��v9@r             g@                           @������@           ��@                           �?WXn�l�@           <�@                           �?�EX@y           �@������������������������       ���Hg[ @�            �v@������������������������       �N-���@�            �n@                           @�0���@@�           p�@������������������������       ��h�ژ�@%           �~@������������������������       �����@v            `h@                           @���.�@           �y@                          �4@V����@             >@������������������������       ��?0-ug�?	             3@������������������������       �?	B0f@             &@                           @�c�lY@�            �w@������������������������       �+�T�Z#@�            �q@������������������������       �P�UYH@C             Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     Ё@      <@      K@     �z@     �Q@     H�@      l@     �@     �u@      @@      ,@     �j@     �t@      3@     �D@     �r@      O@     Py@      g@     w@      n@      ;@      @     �S@     �e@      @      .@      b@      7@     q@     �Q@     @j@     �X@      @      @      O@     �`@      @      &@      \@      *@      m@     �E@     �g@     �R@      �?      @     �J@     �W@      @      @     �R@      $@      `@      ?@     ``@      J@      �?              "@     �C@              @      C@      @     �Y@      (@      N@      7@              @      0@     �D@      @      @     �@@      $@     �D@      <@      3@      8@      @              @      @                      @               @      �?              �?              @      *@      A@      @      @      >@      $@     �C@      ;@      3@      7@      @      @      a@     �c@      (@      :@     `c@     �C@     �`@     @\@     �c@     �a@      4@      @     �X@      `@      (@      1@     @_@      <@     �U@     �X@     @Z@     �\@      2@      �?     �P@     @U@      @      .@     �U@      .@     �J@      Q@     �S@     �I@      *@      @      @@     �E@      @       @     �C@      *@     �@@      >@      :@      P@      @             �B@      <@              "@      >@      &@      G@      .@      K@      :@       @              @      @                      @              ?@      @      2@      @       @              ?@      9@              "@      8@      &@      .@      &@      B@      7@              @     @U@      n@      "@      *@      `@       @     �@      D@     {@     �Z@      @      @      G@      h@       @       @     �T@      @     @@      5@     �u@     �S@      �?              3@      T@      @       @      =@       @     Pq@      @     �d@      ;@      �?              .@      H@               @      1@             @f@       @     �U@      ,@                      @      @@      @              (@       @     �X@      @     @S@      *@      �?      @      ;@     @\@      @      @      K@      @     �k@      0@      g@     �I@              @      $@     �T@      �?      @      @@       @     �f@      $@      a@      @@                      1@      ?@      @      @      6@       @     �E@      @      H@      3@                     �C@     �G@      �?      @     �F@       @      a@      3@     @U@      =@      @               @       @              @                      .@               @      @       @               @       @                                      *@                       @                                              @                       @               @       @       @             �B@     �F@      �?       @     �F@       @     �^@      3@     �T@      9@       @              :@     �A@                      >@      �?     �Y@      (@     �N@      *@       @              &@      $@      �?       @      .@      �?      3@      @      6@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@I£ p~@�	           ��@       	                    �?� +��@d           Ҡ@                           �?~��Y��@�           8�@                            �?m�1�@           x@������������������������       ����1�` @>             W@������������������������       ����E#�@�            Pr@                           @�_��2[@�            `v@������������������������       ���ɱ�@�            `k@������������������������       ����, �?J            `a@
                           �?ƅ��T�@�           �@                           �?��H�g	@@           �~@������������������������       ��}�Lnh@�            �j@������������������������       ����K�
@�            pq@                          �1@L����@H           ��@������������������������       �e�'�@�            �p@������������������������       �a�� �@�           H�@                           @pC���	@g           ��@                           @�E!:s�	@�           ��@                           �?ɿuZ�a	@�           X�@������������������������       ��Ⓗ9"	@�            `w@������������������������       � �"V�@�            Ps@                          �:@���0
@           �{@������������������������       �%7��G�	@�            pq@������������������������       �Za7� �	@f            �d@                            @g�i3@�           ��@                           @駺��V@A           �@������������������������       ���E�c�@6           p~@������������������������       �T、�� @             2@                           @Ȳ	6��@R            �_@������������������������       �x��gF�?)             M@������������������������       ��s/�@)             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �p@     �@      B@     �P@     �{@     �T@     �@     �j@     ��@     �u@     �D@       @      [@     �s@      .@      8@     �h@     �@@     ��@     @W@     p@     �a@      *@             �A@     @T@               @     �K@      @     �u@      3@     �e@      6@      @              ,@     �H@               @      >@      @     @h@      ,@      Q@      $@                              &@              �?      @      �?      F@      �?      8@      @                      ,@      C@              �?      8@      @     �b@      *@      F@      @                      5@      @@                      9@             `c@      @     @Z@      (@      @              2@      7@                      6@             �Q@      @     �Q@      $@                      @      "@                      @             @U@              A@       @      @       @     @R@     �l@      .@      6@      b@      =@     v@     �R@     �t@     @^@      $@       @      B@     �S@      $@      $@     �R@      2@     �Q@     �B@      V@     �K@      @      �?      @     �B@      @      @      <@      @     �E@      4@     �F@      5@              @      =@     �D@      @      @     �G@      .@      <@      1@     �E@      A@      @             �B@      c@      @      (@     @Q@      &@     �q@     �B@     @n@     �P@      @              @     �E@               @      $@             �\@      @     �R@      *@                     �@@     �[@      @      $@     �M@      &@      e@      >@     �d@     �J@      @      2@     `d@     �p@      5@      E@     `n@     �H@     @r@      ^@     �s@      i@      <@      .@     �\@     �e@      0@      B@     �e@      E@     �^@     �W@     �d@     �b@      <@      $@      N@      X@       @      7@     �^@      8@     �U@     �E@     @]@     �T@      $@      @      E@      N@       @      1@      L@      @     �F@      4@     �R@     �A@      "@      @      2@      B@      @      @     �P@      2@     �D@      7@      E@      H@      �?      @      K@     @S@       @      *@     �I@      2@     �B@      J@      H@     @P@      2@      �?      B@      L@      @       @     �A@      @      9@      ?@      <@      ?@      2@      @      2@      5@      @      @      0@      (@      (@      5@      4@      A@              @     �H@     @W@      @      @     @Q@      @      e@      9@      c@     �J@              @     �H@     @U@      @      @      J@      @     �`@      5@      [@     �D@              @      E@     @U@       @      @      G@      @     �`@      4@     �Z@     �D@                      @               @              @      �?              �?      �?                                       @      �?      @      1@             �B@      @      F@      (@                                                      @              ;@              6@       @                               @      �?      @      $@              $@      @      6@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@�e�m�O@�	           ��@       	                    �?�S�f�@�           ��@                           �?tZM9� @           �y@                           �?A�v�w�@H            �[@������������������������       ��W���@              J@������������������������       �.����@(            �M@                           @u���?�            �r@������������������������       ���̖Fc�?z             g@������������������������       ��d�a���?B            �\@
                           @��9; �@�           ؂@                           @}�ᜃ�@�            �w@������������������������       ���)W@F            @]@������������������������       �ؙQ�9@�            Pp@                          �0@H�o�g#@�             l@������������������������       �PI���?             D@������������������������       ���H�9@y             g@                           @R��2�@-           ��@                           �?�����^	@<           ��@                          �<@�|�&{@1           �}@������������������������       �N��8�@           y@������������������������       �A�K	Q�@,            @R@                           �?��lQ�	@           (�@������������������������       ��Wy��h	@
            {@������������������������       ��˵>��	@           Ј@                           �?��΄5�@�           ��@                            @�lAjL@�            0v@������������������������       ��|Z��'@�            �r@������������������������       �B�Qܕf @#            �M@                          �<@i�p�@           h�@������������������������       ���<2o@�           ��@������������������������       ��㓑%a@+             N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     s@     ��@      <@      N@     �z@     @U@     d�@     @i@     ��@     �w@     �@@      @     �N@     �`@       @       @     @U@      @     �y@     �C@     �h@      O@      @              2@      C@               @      @@      �?     �k@      @     @R@      4@                      @      *@               @      5@      �?     �C@      @      0@      "@                       @      @                      "@              6@       @      (@      �?                      @      "@               @      (@      �?      1@       @      @       @                      (@      9@                      &@             �f@      �?     �L@      &@                       @      1@                      �?             @^@      �?      ?@      @                      @       @                      $@             �N@              :@      @              @     �E@     @X@       @      @     �J@      @      h@      A@      _@      E@      @      @      2@     �O@       @       @      E@      �?     �]@      0@     �U@      :@              @      @      .@              �?      $@      �?     �C@      &@      :@       @                      .@      H@       @      �?      @@              T@      @      N@      2@                      9@      A@              @      &@       @     @R@      2@      C@      0@      @               @      &@                                      5@              @      �?                      7@      7@              @      &@       @      J@      2@     �@@      .@      @      0@     �n@      {@      :@      J@     �u@     @T@     ��@     `d@     x�@     �s@      =@      .@     �g@      q@      5@     �C@      l@      O@      o@     �`@     p@     @j@      :@      �?     �L@     �R@       @      *@     �H@      @     �Z@      :@      X@      D@      @      �?      H@      Q@       @      @      D@      @     �Y@      .@     �U@      7@       @              "@      @              @      "@              @      &@      $@      1@      �?      ,@     �`@      i@      3@      :@      f@     �K@     �a@     �Z@      d@     @e@      7@      @     �G@     �U@      "@      @      K@      5@      <@     �E@      J@      R@      "@      $@     �U@     �\@      $@      3@     �^@      A@     �\@      P@     @[@     �X@      ,@      �?      K@     �c@      @      *@      ^@      3@     @x@      >@     �r@     �Z@      @              @     �L@      �?      @      9@      @     `a@      @      X@      5@                      @     �I@      �?              3@      @     �]@      @     �R@      5@                      �?      @              @      @              5@              6@                      �?      H@     @Y@      @      $@     �W@      .@      o@      ;@     �i@     �U@      @      �?      D@     @X@       @      $@      S@      .@     @n@      9@     �h@     �R@      @               @      @       @              3@              @       @      @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJd�;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @p��w>@�	           ��@       	                   �4@��'J�@Y           �@                           �?��r��R@             �@                           �?���]qi@�             q@������������������������       ��p9'Yk@o            @f@������������������������       ��4{4G-@B             X@                           @����5@o           ��@������������������������       �D���@�            0y@������������������������       �Omt\И@s            �g@
                           �?�Up W	@9           ��@                          �:@�`�>�	@w           x�@������������������������       �����)	@�           ȅ@������������������������       ��(̲	@�            `s@                          �5@���>,�@�            Ps@������������������������       ��f�0Or@             I@������������������������       �_��O@�            0p@                           @>�5I�@5           �@                           @�<Z�@�           ܒ@                           �?<*n�	�@�           ��@������������������������       ��
e1��@�            0y@������������������������       �hr���@�             v@                           @�L�V3 @           @|@������������������������       ����Qr�?i             f@������������������������       �td��H @�            0q@                          �=@��u�@M           P�@                          �9@`��(Ԕ@>            @������������������������       ��(�U�@           0z@������������������������       ���X�@-            �S@������������������������       �8�:� `@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        6@     u@     (�@      @@      K@     p}@     @T@     ��@     �g@     `�@     �t@      :@      4@     `n@     �s@      9@     �A@     �u@     �Q@     v@     �b@     `w@      m@      4@      @     �K@     @\@      @      "@     �a@      4@     @h@     �K@      g@     �S@      @              0@      >@                     �B@      @     @U@      &@      R@      3@                      (@      2@                      ?@      @      H@       @      D@      1@                      @      (@                      @             �B@      @      @@       @              @     �C@     �T@      @      "@     @Z@      0@     @[@      F@     @\@      N@      @      @      9@      E@      @      "@      U@      (@     @Q@      9@      U@     �E@               @      ,@     �D@      �?              5@      @      D@      3@      =@      1@      @      ,@     �g@      i@      2@      :@     �i@     �I@     �c@     �W@     �g@     @c@      1@      ,@      b@     @d@      2@      7@     �c@      A@     �Y@     �Q@     �`@     �`@      1@      @     @Y@     ``@      (@      3@     �Z@      2@     �Q@      H@     �[@     �N@      0@      $@     �E@      ?@      @      @      I@      0@     �@@      6@      7@     �Q@      �?              F@     �C@              @      H@      1@      L@      9@     �K@      6@                      @      "@              �?      @      @      @      @      &@                             �D@      >@               @     �D@      $@     �H@      4@      F@      6@               @     �W@     `m@      @      3@     @_@      $@     ��@      D@     `{@     @X@      @       @      P@     @c@      @      @     �T@      @     �@      3@     �r@     �M@       @       @      I@     �V@      @      @     �J@      @     Pr@      2@      g@     �H@       @       @      >@      J@               @      @@      �?     �c@      @     �V@      =@       @              4@     �C@      @      �?      5@      @      a@      (@     �W@      4@                      ,@     �O@              @      >@             �j@      �?     �\@      $@                      @      0@              @      &@             �V@      �?     �H@                               @     �G@                      3@             @_@             �P@      $@                      >@     @T@      @      (@      E@      @     �b@      5@     @a@      C@      @              >@     �S@      @      (@     �B@      @     @b@      5@     ``@      ?@      @              8@      Q@      @      (@      =@      @     �^@      *@     �[@      ?@      @              @      &@                       @      �?      8@       @      5@                                       @      �?              @               @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-��;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�ޏ(�L@�	           ��@       	                    �?L53 1�@}           $�@                           �?\�U��/@�           ��@                          �3@!b�e�@�            �q@������������������������       ��)Ҍ�E@w            �g@������������������������       �m�̛p�@7            �V@                            �?��jϴ	@6           �}@������������������������       ��R�7@W             `@������������������������       �H�o 	@�            �u@
                          �4@��J���@�           h�@                           �?s���?@           ��@������������������������       ��٭8>� @            �z@������������������������       �y�tI@�           @�@                           @�+�03@�            @m@������������������������       �Ն�3"V@@            �Y@������������������������       �w��:��@T            ``@                          �8@���5�@E           ܚ@                          �6@���Z�{@�           �@                           @o�m��V@�            �q@������������������������       ���y� @j            �d@������������������������       ������@N             ^@                            @Q�nL L@8           `~@������������������������       �
CF_ n@�            0u@������������������������       ����D@]            `b@                           @"+�%I	@U           ��@                           @�h�M@�@           @�@������������������������       �pE@;�	@]           ��@������������������������       �gL|�@�            �q@                           �?��?�E�	@G             [@������������������������       ��T$`Q�	@"            �K@������������������������       ���HX�@%            �J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        >@     Pr@      �@      6@     �I@     |@     �R@     X�@      k@     ��@     Pw@      B@      "@     �\@     �r@      (@      :@     �k@      <@     ��@     @Z@     �@      e@      $@      "@      M@     �\@      @      $@     @Z@      .@     �a@      L@     �b@     �V@      @              3@     �F@       @      �?      :@       @     @Q@      4@      Q@      =@                      @      ?@                      6@       @      H@      ,@      F@      6@                      (@      ,@       @      �?      @              5@      @      8@      @              "@     �C@     �Q@      @      "@     �S@      *@      R@      B@     @T@     �N@      @              *@      &@                      6@      �?      3@      2@      ;@      *@      @      "@      :@     �M@      @      "@     �L@      (@     �J@      2@      K@      H@      �?              L@     �f@      @      0@     �]@      *@     X�@     �H@     @v@     �S@      @             �I@      b@      @      (@     �V@      @     �~@      E@     0r@     @Q@                      8@     �E@              �?      7@             �i@      @     @Z@      .@                      ;@     �Y@      @      &@      Q@      @     �q@     �A@     @g@      K@                      @      C@              @      ;@       @     �P@      @     @P@      "@      @               @      .@              @      ,@      @      4@      @      ;@      @      @              @      7@              �?      *@      �?      G@      �?      C@      @      �?      5@     `f@     �n@      $@      9@     @l@      G@     0s@     �[@     �s@     �i@      :@      @     @T@     �^@      @      $@     @X@      (@     �d@      <@     �c@     �S@      $@      @     �A@      I@      @      @      <@      @     �P@      "@     �I@      >@              @      ;@      ?@      �?      @      *@      @      2@      "@     �A@      4@                       @      3@      @              .@      �?      H@              0@      $@              �?      G@     @R@      �?      @     @Q@      @      Y@      3@     �Z@      H@      $@      �?      B@     �G@              @     �E@      @     @R@      0@      S@      <@      @              $@      :@      �?              :@      �?      ;@      @      >@      4@      @      1@     �X@     �^@      @      .@      `@      A@     �a@     �T@      d@     �_@      0@       @      T@      ]@      @      .@     �]@      <@      `@     �Q@      b@     �\@      *@       @     �Q@     @S@      @       @     �V@      7@      L@      L@     @R@      T@      *@              "@     �C@              @      <@      @     @R@      ,@     �Q@      A@              "@      2@      @                      &@      @      (@      *@      0@      *@      @      "@      @      @                      @      @      @      @      @      @      @              *@      @                      @      �?      @      @      (@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJO1�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?0�k�g@�	           ��@       	                    �?��?!	@           ��@                           �?�"�Kפ@v           @�@                          �<@�A�J�@j            �e@������������������������       �[=@�f�@`             c@������������������������       �p�Ͷ��@
             4@                          �:@7q*.^@           �y@������������������������       ��$�+��@�            �u@������������������������       �Չ\k�@,            �N@
                           �?�ԋ�	@�           ��@                          �<@ΰz�]@�            �r@������������������������       �[Ա	�@�            �p@������������������������       �;G�|b@             A@                           @��N� �	@�           H�@������������������������       �ⅷ��	@�           ��@������������������������       �	�O�@
             1@                            �?{
��m@�           �@                           @ �#K�c@&           (�@                           �?��	��@m           (�@������������������������       �g4.l� @�            Pt@������������������������       ��rsU<@�            �@                           �?،q� q@�            Pr@������������������������       ��Ļ9�@_            �b@������������������������       �VV �y@Z             b@                          �3@�����`@�           �@                           �?���@            �y@������������������������       ���I��?a             c@������������������������       ��5��6T@�            @p@                           @J�q�ڀ@�           0�@������������������������       �[7[)J	@_           ��@������������������������       �t[�~(;@,            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     ��@      8@      L@     0{@     @V@     ��@     `m@     ȉ@     0w@      C@      0@     �c@     �l@      (@      ?@     `l@      J@     `k@     @b@     0r@      h@      :@      @      D@     �T@      @      $@     �S@      @     �]@     �F@     @_@      Q@      @              .@      6@                      .@              H@      "@     �H@      *@      �?              &@      2@                      &@             �F@      "@      H@      "@      �?              @      @                      @              @              �?      @              @      9@      N@      @      $@     �O@      @     �Q@      B@      S@     �K@      @       @      7@     �L@       @      $@      I@      @     �P@      <@      Q@      C@      @      @       @      @       @              *@      �?      @       @       @      1@              &@     @]@     @b@       @      5@     �b@      H@     @Y@     @Y@     �d@      _@      5@             �@@     �L@       @      @      E@      �?     �G@      3@     �O@      :@      @             �@@      J@       @      @      A@      �?      G@      .@      N@      0@      @                      @              @       @              �?      @      @      $@              &@      U@     @V@      @      ,@     �Z@     �G@      K@     �T@     �Y@     �X@      2@      @     �T@     @V@      @      ,@     �Z@     �G@     �J@      T@     �X@     @X@      0@      @      �?                                              �?       @      @      �?       @      �?      b@     �r@      (@      9@      j@     �B@     �@     @V@     ��@     `f@      (@              R@     `f@      @      0@     @Z@      8@     Pz@     �H@     �r@     @\@      @             �M@     `a@       @      @     @S@      2@     pu@      B@      m@     �S@      @              *@      B@              �?      @      @      d@      @     �T@      .@      @              G@     �Y@       @      @     �Q@      .@     �f@      @@     �b@      P@      @              *@      D@       @      $@      <@      @     �S@      *@     @Q@      A@                      @      6@      �?      $@      .@       @      B@      �?      D@      1@                       @      2@      �?              *@      @      E@      (@      =@      1@              �?     @R@      _@       @      "@     �Y@      *@     �u@      D@      m@     �P@      @              5@      I@              @      <@             �f@      3@     @W@      (@       @              @      $@                       @             @V@      @      C@       @       @              2@      D@              @      :@              W@      *@     �K@      $@              �?      J@     �R@       @      @     �R@      *@      e@      5@     �a@      K@      @      �?      D@      P@      @      @      P@      &@     `c@      2@     �_@     �J@                      (@      $@      �?              &@       @      ,@      @      *@      �?      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Z����a@�	           ��@       	                     �?czsU�@s           T�@                          �3@;h�]o@�           ��@                           �?X�:@�@�            �k@������������������������       �}h���@,            �Q@������������������������       �����@]            �b@                           �?���Q	@           0}@������������������������       ���IC��@T            �`@������������������������       �t��=;�	@�            �t@
                          �1@j�G��@�           �@                          �0@�4�F��@l            �e@������������������������       �!�r��|@"            �M@������������������������       ��Uvv��@J            �\@                          �;@�� �F	@`           0�@������������������������       �����+�@�           Б@������������������������       �]?���z	@�             k@                          �4@>���d@6           |�@                          �1@�nNޅ�@]           ��@                           @5y�?�             v@������������������������       �ك����?w             e@������������������������       �~�'�?r            �f@                           �?�5_��@t           ��@������������������������       ��^_WoD@�            �t@������������������������       ��5�,@�            �p@                           @��AO�@�           `�@                           �?i[�*@�           ��@������������������������       �Y�C ES@�            �m@������������������������       ��Q�J0*@           `z@                           !@f����	@0            �U@������������������������       ����m��@)             S@������������������������       � ۉ����?             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �p@     ��@     �D@     �F@     �}@     @W@     �@     �m@     X�@     u@     �B@      ,@     @i@     �s@      <@      A@     0t@     @P@      x@     @i@     `w@      n@      @@      @      K@     @Z@      @      "@     �W@      2@     �`@     �R@      _@      K@      0@              "@      ?@                      >@             �K@      =@      L@       @      @               @      @                      ,@              2@      @      8@       @                      @      ;@                      0@             �B@      6@      @@      @      @      @     �F@     �R@      @      "@      P@      2@     �S@     �F@      Q@      G@      (@      �?      (@      9@              �?      *@      �?      D@      �?      @@      @       @      @     �@@     �H@      @       @     �I@      1@     �C@      F@      B@      D@      $@      $@     �b@     �j@      9@      9@     �l@     �G@     �o@      `@     @o@     @g@      0@              *@      7@      �?              1@             �P@      @     �A@      &@                      @      @                      "@              0@      �?      2@      @                      $@      1@      �?               @             �I@      @      1@      @              $@     �`@     �g@      8@      9@     �j@     �G@      g@     �^@     �j@     �e@      0@      @      [@     �c@      2@      0@     �g@      C@     @e@     @[@     �f@     �`@      0@      @      ;@      ?@      @      "@      7@      "@      .@      *@      A@     �E@              �?     @Q@     �n@      *@      &@     �b@      <@     ؃@     �A@     Py@     @X@      @             �@@      a@      @      @      M@      @      {@      *@      k@     �E@                      @     �G@              �?      2@             �g@      @     �R@      $@                      @      4@              �?      "@             �Z@      �?      7@       @                              ;@                      "@              U@      @      J@       @                      ;@     �V@      @      @      D@      @      n@      "@     �a@     �@@                      *@      B@      @       @      :@       @     �a@      "@     �Q@      8@                      ,@      K@      �?       @      ,@      @     �X@             �Q@      "@              �?      B@      [@       @      @     @W@      7@     `i@      6@     �g@      K@      @      �?      9@     �X@      @      @     �R@      2@     @h@      0@     �e@      I@      �?      �?      @     �F@                      0@      *@     �Q@      @     @P@      .@                      3@     �J@      @      @      M@      @     �^@      "@     �[@     �A@      �?              &@      $@      @              3@      @      "@      @      ,@      @      @               @       @      @              2@              "@      @      ,@      @      @              @       @                      �?      @                                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�M�;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@� �B@�	           ��@       	                    @hX"��@T            �@                          �3@2��~ݐ@�           Ԑ@                           �?�=!�V�@�           ��@������������������������       �JP�Ƞ0@�             o@������������������������       �T���@           �{@                            �?0r3z@�             x@������������������������       ��H4wN@E            @]@������������������������       ��MUҬ�@�            �p@
                          �1@q�@�           l�@                           @��A�S @�            �w@������������������������       �x�cP��?�            �o@������������������������       ���)� @I            �^@                          �4@�C�"v@�           �@������������������������       �z���@Y           ȁ@������������������������       �Ϝ'�4@g             e@                            �?K˃��@>           �@                           @��ph(	@?           ��@                           �?kh�p'�	@w           ��@������������������������       ��:�|��@j            �d@������������������������       ���w�
@           �z@                           �?<�Y@�            �r@������������������������       ��~a�4@a            @c@������������������������       ���̽@g            �b@                           @L�7k�@�           Љ@                           �?�'Mʆ@H           H�@������������������������       �愉�K�@R            �^@������������������������       �~|��	@�            �x@                          �;@�ŏ3�@�            s@������������������������       ����� �@�            �k@������������������������       �a%��m@+            �T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     Pt@      �@      7@      M@     Pz@     �U@     ��@     �k@     �@     pw@      =@      @     �`@     �s@       @      5@     �g@      >@     ��@     �W@      �@      g@       @      @     �T@     @b@      @      (@     �`@      8@     @n@      S@     �k@     �]@      @      @     �I@      V@              @     @S@      &@     �e@     �F@     �b@     �T@      �?              5@      >@              �?      :@             �T@       @      N@      5@              @      >@      M@              @     �I@      &@     �V@     �B@     �V@      O@      �?              @@      M@      @      @      M@      *@     @Q@      ?@      R@      B@      @              (@      3@              �?      6@      @      4@      @      5@      &@      �?              4@     �C@      @      @      B@      @     �H@      <@     �I@      9@      @             �I@     �d@       @      "@      L@      @     �{@      2@     `r@     @P@       @              @     �A@              @      4@              g@      @      Z@      2@                      @      ;@              �?      (@             @a@       @      L@      *@                      �?       @              @       @              G@      @      H@      @                      F@     ``@       @      @      B@      @     `p@      *@     �g@     �G@       @              D@      Y@       @      @      8@      �?     �j@      "@     �a@      A@                      @      ?@                      (@      @      I@      @     �G@      *@       @      @     �g@      m@      .@     �B@     �l@     �L@     pt@     �_@     �q@     �g@      5@       @     �[@     �Z@      @      >@      X@     �D@     @b@     �R@      d@      [@      (@       @     @T@      Q@       @      =@     @Q@      @@      O@      P@      X@     �R@      (@              9@      6@              @      "@      �?      >@      *@      E@      2@      �?       @      L@      G@       @      7@      N@      ?@      @@     �I@      K@     �L@      &@              >@     �C@      @      �?      ;@      "@      U@      &@     @P@     �@@                      3@      6@              �?      1@      �?      F@      @      ?@      0@                      &@      1@      @              $@       @      D@       @      A@      1@              @      T@     @_@      "@      @     �`@      0@     �f@      J@     @_@     �T@      "@      @      M@     �W@      @      @     @U@      0@      V@     �D@      O@      L@      "@              ,@      8@                      3@              A@      @      3@      @              @      F@     �Q@      @      @     �P@      0@      K@     �A@     �E@     �H@      "@       @      6@      >@      @       @     �H@             @W@      &@     �O@      ;@               @      2@      6@      �?      �?      4@              S@      @     �J@      6@                      @       @      @      �?      =@              1@      @      $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ2�#IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�;��e@�	           ��@       	                    �?��()�@�           0�@                           @uugo@@           �z@                           @�\�y�@�            �q@������������������������       ��	@�             l@������������������������       ���D�@)            �M@                           �?��A�s @\            �a@������������������������       �L���J�?            �H@������������������������       �� ���� @=             W@
                          �4@}(�<8@�           �@                           @���$�@�             r@������������������������       ��*D�{�@�            @o@������������������������       ���4=,;@             C@                           @�U)]4	@�            0t@������������������������       �z>1��K	@�            �o@������������������������       �=^��M+@.            @Q@                          �1@8���@           z�@                            �?
$���@           P{@                           @&�c��s@i            �d@������������������������       ��z&��/@X             a@������������������������       �[��^ @             <@                           �?�/"��n@�             q@������������������������       ��#_1��@5             V@������������������������       ��?���?{             g@                          �7@���#@�           �@                           �?}��	�%@�           4�@������������������������       �,psn�D@/           �}@������������������������       ��+8V��@�           ��@                           �?K9�h1	@)           ؋@������������������������       �4��s|�@�            �n@������������������������       �8x\G��	@�           8�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �s@     ��@      :@     �S@     �{@     �S@     4�@     �j@     ��@     0w@      :@      @     �W@     �a@      @      1@     @[@      3@     �s@      O@     �e@     @U@      "@       @      A@     @P@              @     �E@      @     @a@      8@      Q@     �B@      @       @      =@     �J@              @      <@      @     @Q@      7@     �A@      ?@      @       @      2@      E@              @      7@      @     �P@      &@      9@      ;@      @              &@      &@                      @      �?      @      (@      $@      @       @              @      (@                      .@             @Q@      �?     �@@      @                              @                       @              ?@              @      @                      @      @                      *@              C@      �?      ;@       @              �?     �N@     �S@      @      (@     �P@      .@     �f@      C@      Z@      H@      @              6@      C@                      8@      �?     �]@      .@      I@      2@      �?              3@      =@                      .@             @\@      .@      E@      0@      �?              @      "@                      "@      �?      @               @       @              �?     �C@      D@      @      (@      E@      ,@     �N@      7@      K@      >@      @      �?     �B@      >@       @      (@      A@      (@      A@      0@     �G@      :@      @               @      $@       @               @       @      ;@      @      @      @              1@      l@      y@      6@     �N@     u@      N@     x�@     �b@     @�@     �q@      1@              "@      F@      �?       @      ?@             �g@      .@     @Z@     �@@      �?              @      2@              @      $@             �P@       @      E@      4@                      @      ,@                       @             �N@      �?      ?@      3@                              @              @       @              @      �?      &@      �?                      @      :@      �?      @      5@              _@      *@     �O@      *@      �?              @       @      �?      @      &@              >@       @      *@      $@                      @      2@                      $@             �W@      @      I@      @      �?      1@     �j@     @v@      5@     �J@      s@      N@     ��@     �`@     �}@     �o@      0@      @     �`@      m@       @      B@     �f@      :@     �w@      P@     pt@      b@      @             �J@      J@              @      >@      @     @e@      ,@     �]@      ;@              @     �T@     �f@       @      >@     �b@      3@     �j@      I@      j@     @]@      @      $@      T@      _@      *@      1@     �_@      A@     @b@     �Q@      c@     @[@      "@              3@      E@              @      =@      �?      M@      "@     �M@      7@              $@     �N@     �T@      *@      *@     @X@     �@@      V@      O@     @W@     �U@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�:��d@z	           ��@       	                    �?|J�,��@W           h�@                          �5@�| ��G	@�           ��@                            �?�Ë�&�@�           ��@������������������������       �a�R5�@�            @l@������������������������       �7]F���@X           ��@                          �:@�V��
@           @�@������������������������       ��T�;�	@D           H�@������������������������       �o�N�	@�            �u@
                           �?F�
�2@c           ��@                           �?��|�)@h             d@������������������������       �)�_�H@;            �X@������������������������       ��3��v�@-             O@                            @C�J�]�@�            `y@������������������������       �q��U,_@�            �r@������������������������       ���.�d@B            �Z@                           �?��̬��@#           T�@                           �?�_]+�; @d           ��@                          �5@5�O�+� @�            0v@������������������������       �t?��FD�?�            @n@������������������������       �;
�f�@F            @\@                           @((�>��?�            �k@������������������������       ��f-���?W             `@������������������������       �/�^��?5             W@                           @�'�B\@�           X�@                           @��DV@�           ȅ@������������������������       ��?�W@�            Pv@������������������������       �6�'u��@�            @u@                            �?ƞ�g^�@           �y@������������������������       �5����K@�             n@������������������������       �=��v&/@p            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �q@     ��@     �B@      K@      }@     �R@     D�@     �m@     h�@     �u@      C@      6@     �i@     Pt@      ;@     �@@      t@     �L@      x@     @i@     �w@     �l@      A@      6@      d@      n@      6@      7@      o@     �H@     �m@     @c@     �q@     @g@      @@      @     @P@     �X@      @      @     �^@      0@      b@     �R@     �e@     �R@      @              7@      <@                      E@       @      A@      6@     �K@      0@      @      @      E@     �Q@      @      @      T@      ,@     �[@     �J@     @]@      M@      @      1@     �W@     �a@      0@      3@     �_@     �@@     �W@     �S@     @\@      \@      9@      @      P@      W@      (@      .@      T@      0@      N@     �F@     �Q@      E@      4@      *@      ?@     �H@      @      @     �G@      1@     �A@      A@      E@     �Q@      @             �G@     @U@      @      $@     @R@       @     `b@      H@     @X@     �F@       @              2@      0@              �?      0@      �?      N@      "@      A@      @                      $@      &@              �?      &@             �C@      @      .@      @                       @      @                      @      �?      5@       @      3@      �?                      =@     @Q@      @      "@     �L@      @     �U@     �C@     �O@     �C@       @              9@      F@      @       @     �H@      @     �G@      >@      K@      >@       @              @      9@       @      �?       @              D@      "@      "@      "@              �?      S@     �i@      $@      5@      b@      1@     x�@      A@     �x@     �]@      @              4@     @T@              @      ;@       @     pr@      @      _@      2@                      (@      K@              @      5@       @     �g@      @      N@      (@                      @     �@@              @      (@             @b@       @      D@       @                       @      5@                      "@       @      E@      �?      4@      $@                       @      ;@                      @             �Z@       @      P@      @                       @      1@                       @             �R@              7@      @                              $@                      @              @@       @     �D@      @              �?      L@     @_@      $@      2@     @]@      .@     �v@      =@     0q@      Y@      @      �?      ;@     �V@      @      1@      T@      &@     �k@      *@     `d@     �P@              �?      0@      A@      @       @      H@      @      `@      @     �U@      9@                      &@      L@      @      .@      @@      @     �W@      @      S@      E@                      =@     �A@      @      �?     �B@      @     @a@      0@      \@     �@@      @              5@      3@      �?      �?      &@      @     �P@      (@     @T@      8@                       @      0@      @              :@      �?     �Q@      @      ?@      "@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJQ� hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�Dŷ@�	           ��@       	                     @��w� @�           ��@                           @�B��@S           ��@                            �?�L�;n�@b           `�@������������������������       ��U���@/           �}@������������������������       �ҭ��
2@3            �T@                            �?Q� /פ@�            �@������������������������       �4OSS�?�            �j@������������������������       �T�S=�@k           X�@
                           @��h�+@6           �@                           �?��}�{m@           �|@������������������������       �_>��@�            `j@������������������������       �ᜁ@�            �o@                           @�����@             E@������������������������       �&����@             <@������������������������       ���h%vO@             ,@                           @�it�I@           H�@                          �:@�*�.>	@"           $�@                           �?|H�˱�@!           ��@������������������������       ��z#�@�           ��@������������������������       ��01¤T@�            �j@                          �<@�q���	@           py@������������������������       ���.�	@k            �e@������������������������       ��\�/��@�            @m@                           @�R>La@�           ؈@                           �?J^%t5@�            �u@������������������������       ��$���@p            `g@������������������������       ��-�}��@f            `d@                          �5@?�:��@            �{@������������������������       ���~2@5            @T@������������������������       ��O8�?@�            �v@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     ��@      <@      C@     �z@     �Q@     �@     �o@     (�@     pv@      <@      @     @Y@     �o@      @      (@     �c@      ,@     @�@      Z@     �v@     @c@       @             @S@     �f@       @      &@     @]@      @     �~@      R@     �p@     @X@      @             �A@     �V@       @      @      T@      @     @_@     �M@     @X@     �K@      @             �@@     @T@       @      @      J@      @      \@     �J@      U@      F@      @               @      $@                      <@              *@      @      *@      &@                      E@     �V@              @     �B@      @      w@      *@     �d@      E@                      @      4@                      "@             �^@       @     �H@      @                     �C@     �Q@              @      <@      @     �n@      &@     �]@     �A@              @      8@     @R@       @      �?     �D@      @     `c@      @@     �Y@     �L@      @       @      8@     �O@       @      �?     �B@      @     �b@      :@     �X@     �I@      �?              .@      =@       @              3@      @     �P@      "@      C@      ;@               @      "@      A@              �?      2@      �?      U@      1@     �N@      8@      �?      @              $@                      @      �?      @      @      @      @      @                      @                      @               @      @      @      @      �?      @              @                              �?       @              �?              @      ,@      h@     Ps@      8@      :@     �p@     �L@     �w@     �b@     `{@     �i@      4@      *@     `b@     �i@      5@      8@      h@      C@     �c@      ^@     �j@      a@      0@      @     @Z@      c@      (@      2@     @b@      6@     �Z@     @R@     @d@     �P@      *@      @      U@     �\@      (@      .@     @\@      ,@     @P@      P@     @_@      G@      (@              5@      C@              @     �@@       @     �D@      "@     �B@      5@      �?       @      E@      K@      "@      @     �G@      0@     �J@     �G@      J@     �Q@      @      @      (@      0@      @      �?      :@      @      A@      0@      6@      <@      �?      �?      >@      C@       @      @      5@      *@      3@      ?@      >@      E@       @      �?     �F@     �Y@      @       @      S@      3@     �k@      <@      l@      Q@      @      �?       @     �J@       @              :@      .@     @[@      *@      Z@      3@              �?      @      ;@                      2@      @     �Q@      @      I@      @                      @      :@       @               @      &@      C@      "@      K@      (@                     �B@     �H@      �?       @      I@      @     �\@      .@      ^@     �H@      @              �?       @              �?      &@      @      *@             �@@      @      @              B@     �D@      �?      �?     �C@      �?     @Y@      .@     �U@      E@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ9�|@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��J��Z@{	           ��@       	                    @��,J@�           ��@                           �?@/§�@�           p�@                           �?:k�@�            Pt@������������������������       �SRƇ/�@8            �X@������������������������       ���H�|�@�            @l@                          �7@��	�f@�            �t@������������������������       �M�����@�             n@������������������������       ��{�_'@9             V@
                            �?����� @Y           ��@                          �6@���J��?M             ^@������������������������       � o>[�?=            �X@������������������������       ��b	�[@             6@                           �?�]t�Ma@           `z@������������������������       ��{�2N@�            `n@������������������������       ������� @q            `f@                            �?2K��|Q@�           :�@                          �5@ �ݍK@�           �@                          �0@S���r@�            �v@������������������������       ��b�@R� @            �C@������������������������       �Q�\!j@�            `t@                           @4��Jp_	@�            @w@������������������������       �߀EѲ	@�            0q@������������������������       �Gǧ�
d@A            @X@                           @��]SU@�           �@                          �?@[B�,��	@�           ��@������������������������       �4��їv	@�           ��@������������������������       �Qo	_�"@             I@                          �:@>C�ۋ/@           ��@������������������������       �
؊zf@�           ��@������������������������       �[�3uӹ@C             [@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     @r@     X�@      7@     �J@     �z@     �U@     �@     �h@     ��@     �v@      E@       @     @U@     @e@      �?      (@      X@      @     �{@      8@     �q@     �P@       @       @     �O@     @Y@              @     @Q@      @     �f@      3@     �b@     �I@      @       @      <@      E@              @     �B@      @      X@      *@     �Q@      :@      �?       @      "@      (@                       @             �@@       @      <@      @                      3@      >@              @      =@      @     �O@      &@     �E@      5@      �?             �A@     �M@              �?      @@       @     �U@      @     @S@      9@      @              :@     �C@              �?      1@             �Q@      @     �P@      1@                      "@      4@                      .@       @      .@       @      &@       @      @              6@     @Q@      �?      @      ;@       @      p@      @      a@      .@      �?                       @      �?              (@      �?     �Q@              9@       @                              @                      @             �P@              2@                                      �?      �?              @      �?      @              @       @                      6@     �N@              @      .@      �?     `g@      @      \@      *@      �?              *@     �C@              @      &@      �?     �\@      �?     �I@      @                      "@      6@                      @              R@      @     �N@      @      �?      :@     �i@     z@      6@     �D@     �t@      T@     P�@     �e@     Ȁ@     �r@      A@      �?     �P@     @Y@      @      "@     @W@      0@      e@     �O@     �^@      T@      &@              2@      I@               @     �K@       @     �Y@      4@     @T@     �@@       @               @      "@                                      0@      �?       @      "@                      0@     �D@               @     �K@       @     �U@      3@     �S@      8@       @      �?     �H@     �I@      @      @      C@      ,@     �P@     �E@      E@     �G@      "@      �?      A@      F@      @      @      =@      &@     �D@      C@      6@     �A@      "@              .@      @      �?              "@      @      9@      @      4@      (@              9@     �a@     �s@      1@      @@     �m@      P@      x@     �[@     �y@      k@      7@      7@     �X@      g@      &@      8@      d@     �J@     �`@     �W@     `f@     �a@      .@      3@     �V@     `f@      "@      8@     �c@      G@     �`@     @W@      e@     �`@      .@      @       @      @       @              �?      @               @      $@      $@               @     �D@     ``@      @       @      S@      &@     �o@      0@     `m@     @R@       @       @      =@     �]@      @      @     �K@      $@     �m@      *@     �j@      N@       @              (@      (@      @      @      5@      �?      1@      @      5@      *@        �t�bub�       hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�"[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?^�v��P@�	           ��@       	                    �?nm縉+@.           ��@                            �?)I�7o�@�           �@                           �?���|5@i            �d@������������������������       �'תz@%            �M@������������������������       ��o��R� @D            �Z@                          �<@Z17�@2           �}@������������������������       ��<�'@            |@������������������������       ��c;b��@             =@
                            �?�9Gi�@�           �@                           @� ���@�            �u@������������������������       ��(_�
@�            �i@������������������������       ���1���?]             b@                           �?�L�nI�@�            `p@������������������������       ��M ,Q@L            �\@������������������������       �D�hJu� @g            �b@                           @�R��P@�           Ƥ@                           @
�5�	@�           ̗@                           �?�����p	@T           �@������������������������       �K_��;�	@N             ^@������������������������       �3Ntj9	@           �@                          �=@�%�U	@v            �f@������������������������       �Y[C%#	@k            @d@������������������������       �"ú�i�@             5@                          �8@Tm;k� @�           ��@                           @2�Y��@I           Ȍ@������������������������       �	���5@�           H�@������������������������       �2�����@�             n@                          �:@-���؂@�            �j@������������������������       �lo� 47@3            @V@������������������������       �5��£�@T            �_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     Ё@      7@     �O@     �{@     @S@     (�@     @k@     x�@     �x@      =@       @     @T@     �g@      �?      &@     �Z@      @     �{@      H@     �r@     @Q@       @       @      B@      Y@      �?      @      K@      �?     @p@      ;@     �\@     �D@               @      @      :@               @      3@      �?     �N@      @     �A@      $@               @      @      *@                      $@              "@      @      ,@      �?                              *@               @      "@      �?      J@              5@      "@                      >@     �R@      �?      @     �A@             �h@      7@     �S@      ?@                      >@     @Q@      �?      @      A@              h@      4@     @S@      5@                              @               @      �?              @      @       @      $@                     �F@     @V@              @     �J@       @      g@      5@     �f@      <@       @              ?@      G@              @     �@@             �V@      $@     �]@      .@       @              =@      <@              @      1@              >@      "@     �R@      *@       @               @      2@                      0@              N@      �?     �F@       @                      ,@     �E@              �?      4@       @     �W@      &@      P@      *@                      "@      <@              �?      *@              =@       @      2@       @                      @      .@                      @       @     @P@      @      G@      @              .@      k@     �w@      6@      J@     �t@     �R@     H�@     @e@     `~@     �t@      ;@      .@     �b@     @l@      3@     �D@      m@     �M@      j@     �a@      i@     �i@      7@      &@     �`@     `h@      3@     �C@     @j@     �G@     @g@     �[@     �g@     �f@      1@      @      1@      $@               @      7@      "@      @      &@      0@      1@      @       @     @]@      g@      3@      ?@     `g@      C@     �f@     �X@     �e@     �d@      ,@      @      1@      ?@               @      7@      (@      7@      @@      &@      6@      @      @      (@      9@               @      6@      @      7@      >@      &@      5@      @              @      @                      �?      @               @              �?      �?             �P@     `c@      @      &@      Y@      .@     �u@      <@     �q@      _@      @              F@     �`@      �?       @     �Q@      &@     s@      $@     `n@     �V@      @              =@     �X@              @      E@      @      n@      "@     �g@      N@      @              .@     �B@      �?      @      <@      @      P@      �?      J@      >@      �?              6@      4@       @      @      >@      @     �C@      2@     �E@      A@                       @      @      �?              (@      �?      3@      1@      5@      *@                      4@      1@      �?      @      2@      @      4@      �?      6@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�y�FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@=��N@�	           ��@       	                    �?���@�           ^�@                           �?Qu���@�           `�@                           �?�l��D@�            @o@������������������������       � �Iy@L            �[@������������������������       ��іm�@S            `a@                          �3@-�I�Q� @T           ��@������������������������       �"/�e @�            `w@������������������������       �J�p=�F@^            �c@
                           @�u?�Ԉ@�           ��@                           �?�KB��@�           І@������������������������       ��C��@L           �@������������������������       ���!��@�            �k@                           �?�4�r
�@�           H�@������������������������       ��E�� l@!            �M@������������������������       �a����@�           p�@                           �?}���@9           h�@                           @aW5��	@3           ��@                           �?7�L�	@�           ��@������������������������       ��p�e@�            @l@������������������������       ��u9M�	@g           ��@                             @�֕ǌQ@9            @V@������������������������       �����,�@%            �L@������������������������       �ǒY���@             @@                           @Km�6��@           �@                           �?����'�@�           @�@������������������������       ������@�             m@������������������������       �?"h�O@j           ��@                           @b<%@             ;@������������������������       �lofON@             &@������������������������       ��1H����?             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@      s@     8�@      :@     �I@     �{@      V@     ��@     @l@     H�@     Pv@      9@      $@     @^@      u@      &@      4@     �j@      <@     H�@     �V@     �~@      f@      "@              H@      Z@      �?      "@     �N@      @     Pt@      2@      f@      @@                      ;@     �@@      �?      @      ?@      �?     �N@      ,@     �M@      1@                       @      &@      �?      @      .@      �?      :@      $@      9@      $@                      3@      6@               @      0@             �A@      @      A@      @                      5@     �Q@              @      >@      @     �p@      @     �]@      .@                      .@      E@              @      0@             �g@      @     �W@      (@                      @      =@                      ,@      @     �R@      �?      8@      @              $@     @R@     @m@      $@      &@     �b@      7@     @x@      R@     �s@      b@      "@      $@     �F@      \@      @      @     @Y@      1@     `b@     �N@     �_@     @W@      @      $@     �A@     �Q@      @      @     �T@      ,@     @T@      D@     �V@     @Q@      @              $@     �D@      �?       @      2@      @     �P@      5@     �B@      8@                      <@     �^@      @      @      I@      @      n@      &@     �g@      J@      @               @      .@                      @      @      "@      @      4@                              :@     �Z@      @      @      F@       @      m@       @     @e@      J@      @      (@      g@     �n@      .@      ?@     �l@      N@     �r@      a@     �q@     �f@      0@      (@     @Z@     �`@      *@      3@     �`@     �E@     @V@     @W@     �]@     �\@      ,@      "@     �X@     �\@      (@      3@     �]@     �C@     �T@      Q@     �\@     @[@      (@              =@     �A@      �?      @      =@      @      3@      ,@      G@      B@      @      "@     @Q@      T@      &@      ,@     �V@     �@@      P@      K@     @Q@     @R@      @      @      @      4@      �?              *@      @      @      9@      @      @       @              @      &@      �?               @      @       @      4@       @      �?       @      @      �?      "@                      @              @      @      �?      @                      T@     �[@       @      (@     @X@      1@      j@     �E@     �d@     �P@       @             �P@     �Z@      �?      (@     �W@      1@      j@     �C@     @d@     �P@       @              (@      <@                      6@      @     @W@      "@     �H@      .@                     �K@     �S@      �?      (@     @R@      (@      ]@      >@     @\@     �I@       @              *@      @      �?               @                      @      @                              �?       @      �?              �?                      @      @                              (@       @                      �?                      �?                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�^�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�0j�*S@�	           ��@       	                    �?Nx�*��@�           ��@                          �<@hZ@�@�           P�@                           �?�2I��.@�           ؂@������������������������       �Rf�:,�@           {@������������������������       ��R7|F@j            @e@                           �?���,�@2            �S@������������������������       �˞2�@             C@������������������������       ��%@�h�@            �D@
                          �9@o���_	@�           ��@                           �?wo��h�@           �@������������������������       ���I0	@%           ��@������������������������       �z�I9�@�            pv@                           @lA*e
@�            �v@������������������������       ��E��&�@9            �T@������������������������       �����=�	@�            `q@                           @^�1�S�@-           �@                           �?D���ԅ@�           ,�@                            �?����N5�?�            `x@������������������������       ��1��B��?9             V@������������������������       �t<`��P�?�            �r@                           @9%i}�@�           (�@������������������������       �B�ь2@�           ��@������������������������       �'S�@             5@                          �5@�G��9@F            @                           �?�2`�v@�            `p@������������������������       ���2��@X            �`@������������������������       ���H� w@Z            �_@                          �=@���2@�            @m@������������������������       �M����@�            �j@������������������������       ���e#��@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@      �@      9@      M@     0|@      U@     ��@     �k@     ؈@     �w@      =@      3@     �l@     pt@      .@      G@     �s@      N@     �x@     �g@     Pw@     p@      ;@       @      R@      X@              @      S@       @     �e@     �B@      a@     @Q@      @       @     �P@      V@              @     �O@       @     �d@      ;@     @`@     �F@      @       @     �I@     �Q@              @      H@      @      Y@      9@      V@     �A@      @              0@      1@                      .@      @     @P@       @      E@      $@                      @       @              @      *@               @      $@      @      8@      �?              �?      @               @      @               @      @      @      ,@                      @      �?              �?       @              @      @      @      $@      �?      1@     �c@     �l@      .@     �C@     �m@      J@     �k@      c@     �m@     �g@      6@      @      Z@     �g@      "@      <@     �h@      >@      h@     �Z@      i@     �`@      1@      @     �T@     �[@      @      :@     `b@      8@      `@     �Q@     �`@     �X@      1@              5@     @S@       @       @      I@      @      P@     �B@     �P@      A@              (@     �K@     �E@      @      &@      E@      6@      >@     �F@     �A@     �K@      @      @      .@      0@       @       @      $@      @              (@      &@       @      @      "@      D@      ;@      @      "@      @@      .@      >@     �@@      8@     �J@       @             �P@      k@      $@      (@      a@      8@     0�@     �@@     `z@     �^@       @              D@     `c@              @     @V@      ,@     �}@      1@     0r@     �R@      �?              *@     �G@                      2@      @      k@      @      S@      $@                              &@                      @             �L@              @       @                      *@      B@                      *@      @      d@      @     @Q@       @                      ;@      [@              @     �Q@      $@     `p@      (@     �j@      P@      �?              ;@      [@              @      Q@      @      p@      &@     `j@     �N@      �?                                              @      @      @      �?      @      @                      :@      O@      $@      "@     �G@      $@     �`@      0@     ``@     �H@      �?              $@      @@      @      @      5@       @     �X@      @     �O@      2@      �?              @      (@      @      @      ,@              I@       @     �B@      $@                      @      4@               @      @       @     �H@      @      :@       @      �?              0@      >@      @      @      :@       @      B@      "@      Q@      ?@                      (@      <@      @      @      9@      @      B@      "@     �P@      6@                      @       @       @              �?      �?                       @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ[ hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?���K+@�	           ��@       	                   �<@���P�	@           4�@                           �?ȢH`ڼ@�           ��@                           �?�`*(z@f           x�@������������������������       ���:�}@�            �l@������������������������       ��4��K�@�            �t@                           �?_�9	5	@           ��@������������������������       �.���lk@�             o@������������������������       �y���T�	@}           ��@
                          �A@�$$��@�            �i@                           @��SR@z             h@������������������������       �qUuk�l@L            �\@������������������������       ���Mv(	@.            �S@������������������������       �B�ޑL��?             *@                           �?��_Ș�@�           ��@                          �2@�7���b@�           (�@                            �?C�r���?�            �q@������������������������       �x��!��?\            @b@������������������������       �߀��S��?Z            �a@                           @ �8��@!           `|@������������������������       �8���ep@N            �^@������������������������       ��o&�@�            �t@                           �?�����@�           \�@                           �?$�`KO�@9            �Y@������������������������       �N��@             B@������������������������       �1j��@&            �P@                           @��ZP*�@�           ��@������������������������       �X�F�t@+           �@������������������������       �	"e�"{@x            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        7@     q@     h�@      4@      L@     0|@     �S@     �@      l@     �@     �w@      :@      6@     �c@     pp@      $@      @@     @o@      H@      l@     `a@     �m@     �j@      3@      0@     �`@     �l@       @      2@     �l@     �D@     �j@     �^@      l@     �c@      2@       @     �@@     @V@      �?      "@     �Z@      @     �[@      D@      W@     �O@      @      �?      *@     �H@              @      N@      @      F@      0@      5@      1@      @      �?      4@      D@      �?      @      G@      @     �P@      8@     �Q@      G@      @      ,@     @Y@     �a@      @      "@     �^@      A@     �Y@     �T@     �`@     @W@      &@             �A@      I@      �?      @     �B@      @     �F@      1@     �@@      7@       @      ,@     �P@     �V@      @      @     @U@      ?@     �L@     @P@     �X@     �Q@      "@      @      7@     �@@       @      ,@      6@      @      *@      1@      (@      L@      �?      �?      7@      ;@       @      ,@      6@      @      *@      0@      (@     �K@      �?      �?      @      2@      �?       @      1@      @      @      @      @     �D@                      1@      "@      �?      @      @      @       @      "@      @      ,@      �?      @              @                                              �?              �?              �?      ]@     `r@      $@      8@      i@      ?@     �@     @U@     ��@     �d@      @              ;@      V@              @     �D@      @     @v@      *@      f@      :@      @              &@      7@              �?      *@             �f@      @     �F@      @      �?              @      ,@              �?      $@              W@              4@       @                      @      "@                      @             �V@      @      9@      @      �?              0@     @P@              @      <@      @     �e@      @     �`@      5@       @              &@      @              �?      "@      �?     �F@      @      C@      @       @              @      M@              @      3@      @      `@      �?     �W@      2@              �?     @V@     �i@      $@      3@      d@      :@     �{@      R@      x@     �a@      @      �?      �?      .@              "@      $@      @      1@      *@      5@      (@              �?               @                      @                      @      ,@      @                      �?      @              "@      @      @      1@      "@      @      @                      V@     �g@      $@      $@     �b@      6@     �z@     �M@     �v@      `@      @             �P@     �e@      "@      $@     @`@      1@     @x@     �G@     �t@      \@                      6@      3@      �?              4@      @      E@      (@     �@@      1@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?iG�t�Y@�	           ��@       	                   �1@9�&;�F@�           �@                           �?�/�G� @�            �p@                          �0@�B�/��@0            �R@������������������������       ���
��@             ;@������������������������       �Y=RzS@            �G@                          �0@�+�(���?v            �g@������������������������       �b6�Xa @(             Q@������������������������       �4@�ۊ5�?N            �^@
                           �?�i��@N           ؍@                            �?���zr@�            v@������������������������       �� ����@I            @]@������������������������       �$�l�L�@�            �m@                           @�~�dC@l           Ђ@������������������������       �g���t@�            Pq@������������������������       �=�����?�            Pt@                          �7@�JqQ@�           
�@                           !@���P@�           �@                          �2@3�/�1@�           ��@������������������������       ��߬}�@�           ��@������������������������       �3 �)	@�           ؒ@������������������������       �����
�?
             2@                           @.�~|<�	@           P�@                           �?ʐfu��	@\           �@������������������������       ��l3R�@S             a@������������������������       �j����6
@	           @y@                           @\�Q(�+@�            �r@������������������������       ��oF�<@�            `n@������������������������       �{�H5
�@              M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        8@     �s@     ȁ@      >@      D@     `{@      V@     �@     �k@     ��@     �t@     �D@      @     @W@     �d@      @      @     �X@       @     �|@      B@     0q@     �P@      @              @      :@                      7@             �a@      @      F@      .@       @               @      (@                      &@              >@      @      &@      @                      �?      @                       @              "@              @      �?                      �?       @                      @              5@      @      @      @                      @      ,@                      (@             @\@      @     �@@      $@       @                      "@                      @              ?@              ,@      @                      @      @                      @             �T@      @      3@      @       @      @     �U@     �a@      @      @     �R@       @     �s@      >@     �l@      J@      @      @     �I@     �L@      @      @     �D@       @     �K@      3@     �T@     �@@       @      @      (@      0@                      *@              0@      @     �E@       @                     �C@     �D@      @      @      <@       @     �C@      *@     �C@      9@       @              B@      U@      �?       @      A@      @     0p@      &@     �b@      3@      �?              ;@     �B@               @      7@      @     �W@      @      R@      &@      �?              "@     �G@      �?              &@             �d@       @     @S@       @              5@     �k@      y@      8@     �A@     @u@      T@     ��@      g@     (�@     �p@      B@      "@      b@     �r@      2@      9@      k@      D@     �|@      W@     �w@      c@      ,@      "@     �a@     �r@      2@      9@      k@     �@@     �|@      W@     Pw@      c@      (@       @      F@     �W@              @     �O@      @     �i@      :@     �a@      D@       @      @     @X@     �i@      2@      3@      c@      >@     �o@     �P@      m@     @\@      $@              @                                      @                      @               @      (@     �S@     �Y@      @      $@      _@      D@     �Y@     @W@     `a@     @\@      6@      $@      M@     �Q@      @      @     @T@      C@     �G@     �Q@     �M@     �S@      3@      @       @      2@                      @@      @      .@      "@      0@      <@      @      @      I@      J@      @      @     �H@     �A@      @@     �N@     �E@     �I@      ,@       @      4@      @@       @      @     �E@       @      L@      7@      T@      A@      @       @      &@      7@              @     �D@       @     �G@      0@     @P@      @@                      "@      "@       @               @              "@      @      .@       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ9�4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@-���!�@�	           ��@       	                   �1@k
N���@P           ��@                           �?|��r�V@x           ��@                           @޷r!�C@�             q@������������������������       ������+@^            �b@������������������������       ����g���?R            �_@                           �?��ƻ�@�            �r@������������������������       ��*x��S@B            @W@������������������������       �C�C�a�?�             j@
                           @E�G�t�@�           l�@                           �?�@�\a@p           ��@������������������������       �lX�߬	@m           ��@������������������������       ���ᴮ@           �y@                          �4@�?�b�f@h           0�@������������������������       ���6º@           �{@������������������������       �e}��[@N            �a@                           @E�X��@_           ��@                            �?�(R=�	@�           ��@                          �7@VZ/E��	@�            �v@������������������������       �+%�� �@J            @\@������������������������       ��W2
@�            �o@                          �:@���N�	@�           ��@������������������������       ����C�@-           �}@������������������������       ��9�
@�            �q@                           @�m0 _�@�           X�@                            �?��n�[[@           �{@������������������������       �/��Ql@C             \@������������������������       ���4�G8@�            �t@                            �?���:Q@�             j@������������������������       �|�gV?@@            @Y@������������������������       ��O/*m@@             [@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@     `s@     8�@     �C@     �H@     P{@     �W@     `�@      k@     X�@     �w@      >@      @     @]@      s@      ,@      6@      j@     �D@     Є@      W@     �~@     `d@      $@              8@     �R@       @      �?     �A@      �?     �n@      5@      b@      <@                      $@     �D@       @              3@      �?     @_@      (@      K@      $@                      "@      8@       @              &@      �?     �N@      (@      4@       @                      �?      1@                       @              P@              A@       @                      ,@      A@              �?      0@             �]@      "@     �V@      2@                      &@      (@              �?      "@              7@      @      8@      "@                      @      6@                      @              X@      @     �P@      "@              @     @W@     �l@      (@      5@     �e@      D@     `z@     �Q@     �u@     �`@      $@      @     �R@     �c@      "@      .@     �`@      C@      h@     �P@     �f@     �W@      $@      @     �K@     �Q@      @      *@     �U@      .@      Y@     �F@     �X@      O@      "@              3@     @V@      @       @      H@      7@      W@      5@      U@      @@      �?              3@     �Q@      @      @     �C@       @     �l@      @     �d@     �D@                      0@      I@      @      @      9@             �g@      @     �\@      A@                      @      4@              �?      ,@       @     �D@      �?     �J@      @              5@      h@     �n@      9@      ;@     �l@      K@      s@      _@     �s@     �j@      4@      4@     @b@     `c@      1@      5@      d@      D@      ^@     �X@     @f@     �b@      1@      @      D@      F@      @      "@     �I@      .@     �G@      C@     �P@      E@      @      �?      1@      *@              �?      6@              5@      (@      0@      $@              @      7@      ?@      @       @      =@      .@      :@      :@      I@      @@      @      0@     �Z@     �[@      *@      (@     �[@      9@     @R@     �N@      \@      [@      $@      �?     �R@     �U@      @      @     �P@      0@     �G@     �B@     �R@      J@      @      .@      ?@      9@      @      @      F@      "@      :@      8@     �B@      L@      @      �?     �G@      W@       @      @     �P@      ,@     @g@      9@     `a@     �O@      @      �?      2@     @P@      @      @      D@      ,@      c@      1@     @W@     �A@                      @      2@       @              .@      @      G@      @      $@      "@              �?      .@     �G@      �?      @      9@       @     �Z@      ,@     �T@      :@                      =@      ;@      @       @      ;@              A@       @      G@      <@      @              3@      &@       @              $@              @      @      B@      0@                      $@      0@      @       @      1@              >@      @      $@      (@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�L	h8@�	           ��@       	                   �1@�p%�@a           *�@                           �?���Ys�@�            �s@                           @��ڌ��@O             `@������������������������       �����+�@$             L@������������������������       �2�F��@+             R@                           �?x.����@h             g@������������������������       �q�/��K@             N@������������������������       �Ą���@L             _@
                           �?�j��0*	@�           t�@                          �;@������	@z           (�@������������������������       ��*� 	@�           (�@������������������������       �*yQ�
@�             p@                           @��.�3;@0           0}@������������������������       �����/B@�            Pr@������������������������       �
V����@p            �e@                          �6@���f�@*           К@                           @��ሑY@           P�@                          �1@/D���� @"           �@������������������������       �JY8���?�             q@������������������������       �d��0�@z           ��@                            @��bT�@�            u@������������������������       �'m�_n�@�            @p@������������������������       ���W�� @5            @S@                          �<@�V�&�@)            ~@                            �?l�43�@�            �x@������������������������       �ȂRw|�@7            �V@������������������������       �n��s�@�             s@                            �?��")Dv@4             U@������������������������       ���7Tc@             D@������������������������       �O��j�@             F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @t@     ��@      <@     �E@     �{@      S@     �@     �j@     `�@     �u@     �A@      5@      l@     �t@      3@      @@     `r@      N@     x@     �e@     0w@     �o@      =@      �?      ,@      I@                      B@      �?     �X@      1@     �O@      ?@              �?      @      6@                      4@      �?     �B@      &@      1@      .@                               @                      &@              4@      "@      @       @              �?      @      ,@                      "@      �?      1@       @      &@      *@                      $@      <@                      0@              O@      @      G@      0@                      @      @                       @              2@      @      2@      $@                      @      7@                      ,@              F@      @      <@      @              4@     `j@     �q@      3@      @@      p@     �M@     �q@     �c@     @s@     �k@      =@      4@     �d@     �i@      2@      >@     @h@     �G@     `f@     @\@      m@     @g@      :@      &@      a@     `e@       @      4@     �d@      @@     `d@      W@      j@     �`@      6@      "@      >@     �A@      $@      $@      >@      .@      0@      5@      8@      J@      @              F@      S@      �?       @      P@      (@     �Z@     �F@      S@     �B@      @              4@     �F@                      H@      "@     @S@      .@      J@      9@       @              8@      ?@      �?       @      0@      @      >@      >@      8@      (@      �?             �X@      n@      "@      &@     �b@      0@     0�@     �B@     �y@     �W@      @              M@     `f@      @      @     �T@      "@     ��@      1@     �r@     �E@      @              E@     @`@       @             �G@      @     �y@      @      l@      <@      �?              (@      :@                      "@             �c@             �M@      "@                      >@      Z@       @              C@      @     p@      @     �d@      3@      �?              0@     �H@      @      @     �A@      @     �^@      (@      R@      .@      @              (@      E@       @      @      @@      @      U@      (@     �J@      &@      @              @      @       @              @              C@              3@      @                     �D@     �N@      @      @     �P@      @     �[@      4@     @\@     �I@       @              A@      L@       @      @      D@      @     �V@      4@     �X@     �D@       @               @      @      �?              (@      @      6@              7@      0@                      :@     �I@      �?      @      <@      @      Q@      4@      S@      9@       @              @      @      �?              ;@              4@              ,@      $@                      @      @                      .@              @              $@      @                      @      �?      �?              (@              .@              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ(��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�RwS@�	           ��@       	                     @+��1��@C           ��@                           �?����@�           |�@                            �?���V��@W           8�@������������������������       ���@[/ @w             i@������������������������       �	*̃��@�            �u@                           @���[+�@�           ��@������������������������       ��D����@{           (�@������������������������       �÷� >@             3@
                           �?X类��@c           0�@                          �1@�
K�@q             f@������������������������       ��h�Ӂ?@            �F@������������������������       �P͠��@T            �`@                          �2@�n���@�            Pw@������������������������       ��'р��@w             f@������������������������       �T��]	@{            �h@                          �<@*�@o��@Y           �@                           �?���=V@}           ��@                           �?c��	�@�            Px@������������������������       ���
�_@w            �f@������������������������       �����I�@�            �i@                           @y�L�@�           x�@������������������������       �� #��@%           Ћ@������������������������       ����{��@a            �d@                            �?����>�@�            v@                           @�ZGʫ�@~            @j@������������������������       �/w7��@?             [@������������������������       ��k+�Es@?            �Y@                           @F���c@^            �a@������������������������       �]��qD�@L            @\@������������������������       �� k@             >@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@      t@     ~@      D@     �J@     }@     @R@     �@     �l@     8�@     �w@      ;@      @     �\@     @q@      .@      7@      k@      8@     Ȅ@     �V@     �@      d@      (@      �?      V@     �i@       @      ,@     @b@      *@     `�@     �O@     �w@      ]@      "@              <@      O@               @     �B@      �?     �l@      .@     �`@     �D@       @              @      7@                      @             �V@      �?      L@      2@                      8@     �C@               @      >@      �?      a@      ,@     �S@      7@       @      �?      N@     �a@       @      (@     @[@      (@     �r@      H@     �n@     �R@      @             �M@     �a@       @      &@     @Z@      "@     Pr@     �G@     �n@     �Q@      @      �?      �?                      �?      @      @      @      �?      �?      @              @      :@     �Q@      @      "@     �Q@      &@     �a@      <@     �`@      F@      @              $@      6@              @      .@              P@       @      E@      *@                       @      @                       @              5@      @      @                               @      3@              @      @             �E@      @      B@      *@              @      0@     �H@      @      @      L@      &@     @S@      4@      W@      ?@      @               @      9@       @       @      9@              G@      @     �H@      *@              @       @      8@      @      @      ?@      &@      ?@      ,@     �E@      2@      @      "@     �i@     �i@      9@      >@      o@     �H@     �t@     �a@     Pt@      k@      .@      "@      d@      d@      3@      5@     �h@     �C@     pr@      Z@     �q@     `a@      (@      �?      E@      E@       @      �?     �G@      "@     @Z@      &@      Y@      :@      @      �?      =@      3@      �?      �?      C@      @      :@      "@     �C@      ,@      @              *@      7@      �?              "@      @     �S@       @     �N@      (@               @     �]@     �]@      1@      4@     �b@      >@     �g@     @W@     `g@     @\@      "@       @     �W@     �W@      ,@      4@     �_@      6@     @e@      Q@      e@     @X@      @              7@      7@      @              8@       @      4@      9@      3@      0@      @              G@     �F@      @      "@      I@      $@     �@@      B@      C@     @S@      @              9@      <@              @      3@      @      ,@      9@      9@      M@      @              $@      ,@              @      @       @       @      ,@      @      C@       @              .@      ,@                      (@      @      @      &@      2@      4@      �?              5@      1@      @      @      ?@      @      3@      &@      *@      3@                      4@      1@      @      @      9@      @      (@      &@      @      ,@                      �?              @              @              @               @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��__hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@U]<�TE@�	           ��@       	                    �?���q��@�           ��@                          �3@����@�           (�@                           @b�i���@2            ~@������������������������       ��c�oh�@�            `x@������������������������       � a48/@9            �V@                           @^G`G�@T            �`@������������������������       �D5�f@5             T@������������������������       ��֤�@            �J@
                           �?^W��e@           �@                            �? $K0�} @           `|@������������������������       �3����V�?Q            �_@������������������������       ���l�� @�            �t@                            �?��J0T@�            �@������������������������       �٤e��@           P|@������������������������       ��׫�@�            �s@                           �?��٥&�@            <�@                          �7@+�;�@v           ��@                           �?�{S�@�            �o@������������������������       �'i:�F@T             a@������������������������       �DjF{P@J             ]@                           �?@4W0@�            Pu@������������������������       �V�;e>*@p            �f@������������������������       ��ӓ��@h            �c@                          �<@_�A�pT	@�           0�@                           �?މ��	@           ��@������������������������       ��a����	@;            �W@������������������������       ���8��@�           �@                           �?�)}&H	@�            �m@������������������������       ���t��@,             R@������������������������       ��i`�N	@h            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      r@     p�@      8@      M@     0|@      U@     Џ@     �k@     ��@     Pw@      >@      �?     @[@      l@      @      &@     �f@      3@     ��@      S@     �x@     @a@      "@      �?      N@     �P@      @      @     �X@      (@     �`@      K@     �Y@     @Q@      "@      �?      B@      J@      @      @     �S@      &@      ^@      B@     �Q@     �O@      @      �?      ;@      B@       @       @     @P@      $@     �X@      ;@     �P@      K@                      "@      0@       @      �?      *@      �?      5@      "@      @      "@      @              8@      ,@                      5@      �?      ,@      2@      @@      @      @              0@      *@                      (@      �?      $@       @      2@      @      @               @      �?                      "@              @      0@      ,@      �?                     �H@     �c@      @       @     �T@      @     p�@      6@     �r@     @Q@                      3@      J@               @      7@             �k@      @     �[@      4@                      @      0@              �?      @              M@              C@      @                      0@      B@              �?      4@             �d@      @     @R@      *@                      >@     �Z@      @      @     �M@      @     �r@      2@     @g@     �H@                      ,@      L@      @       @     �E@      �?     �f@      $@     @\@      =@                      0@     �I@              @      0@      @     @^@       @     @R@      4@              0@     �f@     �t@      1@     �G@     �p@     @P@     `v@      b@     `x@     `m@      5@      @     �D@     �Y@      �?      "@     �P@      @     �b@      8@     �a@     �H@      �?              2@     �K@      �?      �?      0@      @     �T@      �?      N@      0@                      @     �@@              �?      (@      @     �L@              5@      @                      .@      6@      �?              @              9@      �?     �C@      "@              @      7@     �G@               @     �I@      @     �P@      7@     �T@     �@@      �?      @      2@      ?@               @     �B@      �?      6@      ,@      <@      4@      �?              @      0@                      ,@       @      F@      "@     �K@      *@              *@     �a@     �l@      0@      C@     `i@     �M@     @j@     @^@     �n@     @g@      4@      (@      [@     �h@      .@      ;@     @d@     �E@     `h@     �X@     `l@     �b@      1@      @      2@      "@               @      *@      @       @      (@      &@      $@       @      @     �V@     `g@      .@      9@     �b@      C@     `g@     �U@      k@     @a@      .@      �?      @@     �A@      �?      &@     �D@      0@      .@      7@      4@      C@      @      �?      (@      .@      �?              *@      "@       @      @      @      "@                      4@      4@              &@      <@      @      *@      2@      .@      =@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ*62hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @'G��uM@�	           ��@       	                    @$�$�@�           ڥ@                           �?������@�           z�@                           @(�^�	@>           ��@������������������������       �����?4@r           ��@������������������������       �lR9_��	@�            0t@                           @�d�?�@�           ��@������������������������       �d���@
           z@������������������������       �����@{           �@
                           �?�n����@             H@������������������������       �^�z|�X�?             (@                           @�Jv@             B@������������������������       �<K)= @             9@������������������������       ���^~@             &@                          �9@%��@�           p�@                           �?U;�@2           H�@                          �0@B���=|@�             q@������������������������       ��F��h��?             4@������������������������       �@D~�?�@�            �o@                           �?n$|�@~           ��@������������������������       �����	�@�            @n@������������������������       ���[��@�            Pv@                          �<@����
@�            `n@                           @ǿ?9u�@T            �`@������������������������       �hu2�@A            �Y@������������������������       �p?Ǌ�.@             ?@                           @j��uxn	@E            @[@������������������������       �Dj��oF	@3             T@������������������������       � �����@             =@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     @s@     x�@      B@      H@     �}@      T@     ��@      k@     ��@     �t@     �C@       @     `k@     �w@      6@      ;@      t@      O@     ��@     �a@     ��@     �l@      8@       @     �i@     �w@      6@      ;@     �s@     �M@     ��@     �`@     ��@     �l@      2@      @     �W@     @b@      .@      (@     `a@      =@      a@     @R@     �a@     �[@      .@      @     �M@     �W@      @       @      W@      7@     @X@      =@     �[@     @R@      @      @     �A@     �I@      (@      @     �G@      @     �C@      F@     �@@      C@      &@      �?      \@      m@      @      .@     `f@      >@     H�@      N@     p|@     @]@      @              >@      E@              @      J@      ,@     �[@      ?@     �W@     �A@       @      �?     �T@     �g@      @      "@     �_@      0@     �@      =@     �v@     �T@      �?              *@                              @      @      @      "@       @      �?      @                                               @       @      �?              �?              @              *@                               @      �?      @      "@      @      �?                      "@                                              @      @      @      �?                      @                               @      �?               @       @                       @     @V@     �b@      ,@      5@      c@      2@      p@     �R@     �j@     �Z@      .@      @      O@     @`@      "@      &@      `@      $@     �j@     �E@     @g@     �P@      @              2@      >@      �?      @      6@              Y@      "@      S@      .@                                                      @              &@      �?      @                              2@      >@      �?      @      2@             @V@       @      R@      .@              @      F@      Y@       @       @     �Z@      $@     �\@      A@     �[@     �I@      @      @      *@     �D@      @      @      F@      @      G@      $@     �H@      6@       @       @      ?@     �M@       @      @     �O@      @     @Q@      8@     �N@      =@      @      @      ;@      2@      @      $@      7@       @     �D@      @@      <@      D@       @              *@      @      @       @      (@      @     �A@      *@      .@      7@       @              *@      @      �?              $@      @      2@      &@      (@      4@       @                               @       @       @              1@       @      @      @              @      ,@      ,@       @       @      &@       @      @      3@      *@      1@              @      $@      @       @       @      $@       @       @      1@      @      (@                      @      @                      �?              @       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJۇ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@3�S`�Q@�	           ��@       	                    �?���;�@S           �@                           @{�T��@�            �@                           �?�Ǡ���@            }@������������������������       �7�<�Z@�            �k@������������������������       ����� L@�            �n@                          �2@7��}&�?�             s@������������������������       �8��b��?v            @g@������������������������       ��b<S�F�?H             ^@
                           @�D�t�@v           �@                            �?�imn��@�           `�@������������������������       ��eQ�.@�            �j@������������������������       �ĻN�@E           ��@                           @��eX�s@�           ��@������������������������       �������@m            �f@������������������������       �$�.v��@=            ~@                           @r�Ŷ�@H           �@                           �?ǵ���N@�           �@                          �<@�ىQ@2           �}@������������������������       ��0��ٍ@�            �w@������������������������       �c��d�J@>            @W@                            �?6�Y��@�           ��@������������������������       ����N$7	@�            �r@������������������������       �-�"���@�           ؇@                           �?�,���	@q            �g@                           �?m�H27�@/            �S@������������������������       �����@             5@������������������������       ��9��*�@"            �L@                            �?��w8]@B            �[@������������������������       ���MO�s@             7@������������������������       ���q�J�@4            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     ��@      :@     �J@     �|@      R@      �@     `l@     Ј@     �w@      >@      $@     @[@     pt@       @      7@     �j@      ?@      �@     �X@     0~@     `d@      *@             �C@     @]@              @      K@      @     �t@      6@     `d@      D@                     �@@     �S@              @      D@      @     �c@      3@     �Y@      =@                      .@      D@              @      9@      @      S@      *@     �@@      *@                      2@     �C@              �?      .@              T@      @     @Q@      0@                      @      C@              �?      ,@             �e@      @     �N@      &@                      @      ,@              �?      *@              [@      @     �A@      @                      �?      8@                      �?              P@              :@      @              $@     �Q@     @j@       @      2@      d@      ;@     �w@      S@      t@     �^@      *@      $@     �G@     @\@      @      .@     @]@      2@      b@     �P@     �_@     @S@      "@              1@      5@              �?     �C@      @     �D@      6@      D@      8@      �?      $@      >@      W@      @      ,@     �S@      (@     �Y@     �F@     �U@     �J@       @              7@     @X@      @      @      F@      "@      m@      "@     @h@      G@      @              "@     �B@                      @      @      M@      @     �E@      ,@      @              ,@      N@      @      @      C@      @     �e@      @     �b@      @@              (@     �g@     @m@      2@      >@     `n@     �D@      r@      `@     ps@      k@      1@      @      d@     �i@      *@      >@      j@     �A@     �p@      Y@     �r@     `i@      *@      �?      D@     �S@              @     �K@      @      Z@      2@      \@     �K@      @      �?     �@@      P@               @     �E@      @     �V@      $@     @Y@      @@      �?              @      ,@              �?      (@      �?      ,@       @      &@      7@       @      @     @^@     �_@      *@      ;@     @c@      =@     @d@     �T@     �g@     �b@      $@       @      C@     �D@      @      @     �A@      (@      M@      <@      B@     �C@      @      @     �T@     @U@      $@      4@     �]@      1@      Z@      K@      c@     @[@      @      @      <@      >@      @              A@      @      6@      =@      $@      ,@      @      @      @      4@      �?              "@       @       @      .@               @      @      �?       @       @      �?              @      �?              @               @              @      @      2@                      @      �?       @       @              @      @              7@      $@      @              9@      @      ,@      ,@      $@      @                      @              @                      �?       @      @      @      @                      3@      $@      �?              9@      @      (@      $@      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�p;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@?>��6@�	           ��@       	                    �?�6���@�           ��@                          �2@JМ>ʶ@P           ��@                            @�"Ec� @           �z@������������������������       ���� @�            ps@������������������������       �$34s'�@H            �\@                           @&�,�a@I            �[@������������������������       ��g���@/             R@������������������������       ���u/AC�?             C@
                           @��W�@6           ��@                            �?�'f�&�@_           ��@������������������������       ��ԅ7"@�             r@������������������������       �!阽��@�            `q@                           @�Ɠ5j@�            �u@������������������������       ��.�_�@�             m@������������������������       ��5�����?M             ]@                          �8@�k�W8=@           @�@                            @��ұ^�@�           ��@                          �4@Π�C;Q@�           ��@������������������������       �k�ܰ�@�            �q@������������������������       ���!��@           8�@                           �?h�QK�@           �|@������������������������       ���U-@             j@������������������������       ���tO)�@�            �n@                          �:@z��<�@7           ��@                           @:��@X@�            @v@������������������������       ��dyх(	@�             l@������������������������       �
��oA@N            ``@                          �;@d;���@\           p�@������������������������       ��pf�'�@V            `a@������������������������       �f�d=H	@           0x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      r@     ؀@     �A@      J@     �|@     �T@     @�@     @g@     P�@     0w@      ?@       @     @P@     �f@      @      *@     ``@      *@     �@     �M@     Ps@     �\@      @              5@      J@               @      C@      �?     �n@      &@     @`@      @@      �?              *@      C@               @     �@@      �?     �j@      @     �X@      4@      �?               @      8@                      7@             `d@      @     @R@      ,@      �?              @      ,@               @      $@      �?     �H@       @      9@      @                       @      ,@                      @             �A@      @      @@      (@                       @      &@                      @              ,@      @      5@      $@                              @                                      5@      �?      &@       @               @      F@      `@      @      &@     @W@      (@     �r@      H@     `f@     �T@       @       @      @@      U@       @      "@     @Q@      (@      b@     �F@     @V@     �Q@       @      �?      2@      B@       @      @     �A@      @     �T@      2@      E@      E@       @      @      ,@      H@              @      A@      @     �N@      ;@     �G@      <@                      (@     �F@      @       @      8@             �c@      @     �V@      *@                      "@      B@      @      �?      3@             �V@      @     �P@      @                      @      "@              �?      @             @P@              7@      $@              .@     �k@     `v@      >@     �C@     Pt@     @Q@     �~@     �_@     P@      p@      <@      @     �`@     �n@      0@      ?@     �i@     �B@     0w@     �N@     �t@      `@      2@      @      V@     @f@       @      8@     �a@     �A@     �q@      G@     �m@     �R@      @              6@     �E@      �?      @      ?@      @     �V@      *@     �L@      7@              @     �P@     �`@      @      5@     �[@      @@     �g@     �@@     `f@     �I@      @              G@      Q@       @      @      P@       @     @V@      .@      W@      K@      &@              7@      5@       @      @      ;@      �?      H@      @      C@      :@       @              7@     �G@               @     �B@      �?     �D@      &@      K@      <@      @      "@     @V@      \@      ,@       @     �]@      @@     �^@     �P@     �e@      `@      $@              A@     �G@      @      @     �B@      ,@     �H@      @@     �V@      C@      @              @@      D@      @      @      9@       @      4@      =@      B@      5@      @               @      @              �?      (@      @      =@      @      K@      1@              "@     �K@     @P@       @      @     �T@      2@     @R@      A@     �T@     �V@      @      �?      &@      (@                      8@              =@      (@      8@      8@       @       @      F@     �J@       @      @      M@      2@      F@      6@     �M@     �P@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @hl�Y�@�	           ��@       	                    �?rtx�D5@�           Υ@                           @gش�?@J           ��@                          �8@��$�@l           Ȁ@������������������������       ���Y�@           @y@������������������������       ���C4�@T            �`@                          �5@�h���  @�            Pv@������������������������       ��F9��?�            @o@������������������������       ��ĸИ�@A            �Z@
                          �5@K�&�f3@�           ��@                           @D ���@�           t�@������������������������       �,�0��_@�           H�@������������������������       ���n*@�            @y@                           �?}^^Zf	@"           `�@������������������������       ��=��*
@(             O@������������������������       �R�	@�           p�@                           �?���E@�           ��@                          �3@S�/�Q@�             u@                           �?�ˮL
T@Y            �`@������������������������       ��+���@'            �L@������������������������       ��h�Bj�?2             S@                           @rE����@x            `i@������������������������       ��V��k@[             c@������������������������       ���I
�@             I@                          �9@%F�8�@�           ��@                           @^���6!@�           ��@������������������������       �Ж��G�@]           8�@������������������������       ���Wq~@'             L@                           @5��KbL
@t            `f@������������������������       �Gp����@             D@������������������������       ���h�	@Y            `a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     Ps@     ��@      C@     �H@     0~@     @U@     ��@     �k@     ��@     @w@      @@      *@     `j@     0y@      5@      :@     �t@      Q@     H�@     @d@     �@      o@      2@      �?      N@     @_@      @      �?     @V@      @      s@      7@     �k@     �L@       @      �?      J@     �Q@       @      �?      R@      @     @_@      ,@     `a@      J@       @             �D@     �H@       @      �?      I@       @     @\@      $@     �Z@      >@              �?      &@      6@                      6@      @      (@      @     �@@      6@       @               @      K@      �?              1@      �?     `f@      "@     �T@      @                      @     �A@                      "@             �b@      @      F@       @                      �?      3@      �?               @      �?      =@      @     �C@      @              (@     �b@     `q@      2@      9@      n@     �N@     �y@     `a@     0v@      h@      0@       @      Q@     @d@      "@      &@     @\@      8@     �r@      I@     `k@      V@      @              <@      \@      "@      $@     @S@      1@     `e@      :@     �a@      M@               @      D@      I@              �?      B@      @     ``@      8@     �S@      >@      @      $@     �T@      ]@      "@      ,@      `@     �B@     �Z@     @V@      a@      Z@      &@      @       @      @              @      @      @      @      &@      $@      @      �?      @     �R@     �[@      "@       @     �^@     �@@      Z@     �S@     �_@     �X@      $@       @     �X@     `e@      1@      7@      c@      1@     �l@     �M@      j@     �^@      ,@              >@      E@      �?       @      A@             @[@      .@     �Q@      ;@                       @      *@                      @              M@       @     �B@       @                      @       @                      @              ;@       @      &@      @                      @      &@                       @              ?@              :@      �?                      6@      =@      �?       @      ;@             �I@      *@     �@@      3@                      6@      7@      �?      @      5@              >@      &@      5@      2@                              @               @      @              5@       @      (@      �?               @      Q@      `@      0@      .@     �]@      1@     �^@      F@     @a@      X@      ,@      @      F@      Z@       @       @      Y@      $@     �Y@      ?@     �^@      O@      &@      @      C@     �V@       @      @      V@      "@     �X@      :@     �]@      N@      @      �?      @      *@               @      (@      �?      @      @      @       @      @      @      8@      9@       @      @      3@      @      4@      *@      0@      A@      @              @       @      @       @                      �?       @      @      @      @      @      4@      1@      @      @      3@      @      3@      @      (@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�!�IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\�)     C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��,ʤa@�	           ��@       	                   �5@�[벏�@z           �@                           �?V�O%��@�           ��@                           �?���%�,@�            v@������������������������       �U,��@g            �d@������������������������       ��T�@p            @g@                          �1@��X@�           ��@������������������������       ��g�k<@n             f@������������������������       �%��%up@k           `�@
                          �8@_��	��	@�           <�@                           �?O�e�@9           ~@������������������������       �N�}�Te@U            �]@������������������������       �+�{^�=@�            �v@                           �?��k� 
@�           p�@������������������������       �S ,:�i
@D           �@������������������������       �2Q�9�@M            @]@                           �?�S��3@9           ��@                          �4@5��@� @e           ��@                          �0@*&M���?�             u@������������������������       ��jp���?&             N@������������������������       ��Õk3�?�            @q@                          �7@�i�n)@�            `l@������������������������       �jx���h@J            �]@������������������������       �Y�FP^@D            @[@                           @����h@�           (�@                            �?�DA�@8@�           ��@������������������������       ��(@m��@�            `o@������������������������       ��[�r>\@           ��@                           @��l�t@             >@������������������������       �|���7��?             $@������������������������       �;z�0��@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �p@     ؁@     �A@      M@     �|@     �W@     ��@     �k@      �@     �t@      A@      3@     �h@      u@      <@      E@     `t@     @R@     �w@      e@     �w@     @k@      :@      @     �M@     �c@       @      7@     `d@      7@     �n@      U@     �j@      W@      &@              8@      J@       @      @      I@      @      X@      1@     �T@      0@      @              "@      7@       @       @      ;@      @      H@      (@      >@      @      @              .@      =@               @      7@              H@      @      J@      (@              @     �A@     �Z@      @      3@     @\@      1@     �b@     �P@     @`@      S@      @       @      "@      C@      @       @      @      �?     �H@      1@      <@      5@              @      :@     @Q@      @      1@     �Z@      0@     �X@      I@     �Y@     �K@      @      (@      a@     `f@      4@      3@     `d@      I@     �`@     @U@     �d@     �_@      .@      �?     �T@     �U@      @      "@     @U@      (@     �K@      1@      T@     �E@      @              9@      6@      �?              .@              6@       @      8@      @       @      �?     �L@     @P@      @      "@     �Q@      (@     �@@      .@      L@      C@      @      &@     �K@      W@      .@      $@     �S@      C@     �S@      Q@      U@     �T@      $@      &@     �G@     @S@      .@      $@      P@     �@@     �G@     �J@      Q@     �Q@      "@               @      .@                      ,@      @      ?@      .@      0@      (@      �?      �?     @Q@      m@      @      0@     �`@      5@     �@     �J@     �z@     @]@       @              &@     �R@      �?      @      6@      @      r@      .@     �_@      1@       @              @      <@              @      *@             �h@       @     �Q@      @       @                      $@                      @              @@              $@      �?                      @      2@              @      @             �d@       @      N@      @       @              @      G@      �?              "@      @     �V@      @      L@      $@                      @      ;@      �?               @      @      K@      �?      3@       @                       @      3@                      �?              B@      @     �B@       @              �?      M@     �c@      @      (@     @\@      2@     �u@      C@     �r@      Y@      @      �?     �K@     �c@      @      (@      [@      (@     �u@      B@     @r@      Y@      @              5@      =@                      1@      @      X@       @     �J@      7@              �?      A@     �_@      @      (@     �V@       @     �o@      <@     �m@     @S@      @              @      @                      @      @      �?       @      $@                                                              @       @               @       @                              @      @                      �?      @      �?               @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ_qOKhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@ڵ�C�@�	           ��@       	                    �?q(m�@D@�           0�@                          �0@IY~�@           ��@                           �?�Χ��?2             W@������������������������       �#K�e�"�?             J@������������������������       ��}F0�%@             D@                           @���f��@�           ؇@������������������������       ��)L���@            `|@������������������������       ��g�5X�?�            Ps@
                          �1@_�+�=@�           �@                           �?�F�`�@�            �t@������������������������       �M3*�@5            @U@������������������������       ���fF$@�             o@                           �?D?�� �@           Г@������������������������       �4����@=           �@������������������������       �q��!�1@�           ��@                           �?LC�i�@�           Ė@                           @�%����	@�           P�@                           �?{Sz��	@�           ��@������������������������       �<��@�            �m@������������������������       �u����	@           pz@                          �<@��E��@3            �U@������������������������       ��̓�#@%             P@������������������������       �	m��@             7@                           @��q���@�           8�@                            @%��n�@�           ��@������������������������       ����3W�@<           `~@������������������������       �oWiCf@W            `a@                            �?`p��4W@8            �U@������������������������       �V��6@
             2@������������������������       �G�� �@.             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pt@     ��@      9@      O@     0�@      Z@     ��@      h@     ؇@     0v@     �A@      (@     �f@     �t@      (@      B@     pq@      E@     ؇@     @X@     �@      f@      *@             �Q@     �Y@       @      @     �P@      &@     @u@      :@     �g@     �E@                      �?      5@                      @             �F@              $@       @                              .@                       @              =@              @       @                      �?      @                      @              0@              @      @                     @Q@     �T@       @      @     �M@      &@     pr@      :@     `f@     �A@                     �K@     �F@       @      @      G@      &@      `@      3@     �\@      <@                      ,@     �B@                      *@             �d@      @      P@      @              (@     @\@     �l@      $@      ?@     �j@      ?@     pz@     �Q@      t@     �`@      *@              0@     �B@      �?      @      6@      �?     �_@      3@     @T@      :@                      "@       @      �?       @      &@      �?      (@      &@      0@      ,@                      @      =@              �?      &@             �\@       @     @P@      (@              (@     @X@      h@      "@      <@     �g@      >@     �r@      J@     �m@      [@      *@      �?      >@     �T@      @      (@      U@      .@     �[@      (@      \@      I@      �?      &@     �P@     �[@      @      0@     �Z@      .@      g@      D@     �_@      M@      (@      $@      b@     �h@      *@      :@     �m@      O@     �j@      X@     �o@     @f@      6@      "@     �U@     �X@      *@      3@     �b@      C@     �J@     �O@     @W@     �Z@      4@      @     �S@     @V@      *@      3@     �`@      A@      H@     �E@      V@     @W@      ,@      @      7@      >@      �?      �?     �I@      @     �@@      @     �E@     �@@      @      �?     �K@     �M@      (@      2@     �T@      =@      .@     �B@     �F@      N@      "@      @       @      "@                      ,@      @      @      4@      @      *@      @              @      @                      &@      �?      @      4@      @      &@      @      @      @      @                      @      @                       @       @      �?      �?      M@      Y@              @     �V@      8@     @d@     �@@      d@      R@       @      �?     �D@     �T@              @     �T@      7@     �b@      7@      b@     @Q@      �?      �?      >@      N@              @      R@      6@      Z@      .@      ^@     �K@      �?              &@      7@              �?      $@      �?      G@       @      9@      ,@                      1@      1@                      "@      �?      (@      $@      0@      @      �?              @       @                                      @              @      @                      *@      .@                      "@      �?      @      $@      (@              �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�t:hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?GL�G@�	           ��@       	                    �?�8{@           ԓ@                          �7@-����@�            �@                          �5@�r-(�@3           �~@������������������������       �����9�@           @z@������������������������       � �ˬ�8@/            �R@                            @w�@o             f@������������������������       ������@O            @`@������������������������       �%��5@             �G@
                           @p�S�@w           ��@                            �?b>��j]@�            �u@������������������������       �`�f��@u             g@������������������������       �F={M�@g             d@                          �4@\�ݯ� @�            �o@������������������������       ���V�~�?Z            @c@������������������������       ����>�@A            �X@                           @	��U&U@�           ��@                            �?Ȕ;;�d	@�           �@                           @��_�@$           @}@������������������������       �E6� Y@�            �x@������������������������       �4��J/�@)            �Q@                           @�O��	@�           ��@������������������������       ��F���\	@�           4�@������������������������       �=g�q�@            �A@                           @2L�v0C@�           @�@                          �<@�
�R��@           8�@������������������������       �3�Ƙ�@�           ��@������������������������       ��!�p'@             D@                            �?�9=mWz@�            �t@������������������������       �u���l@,            �O@������������������������       ���#&�!@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     0s@     H�@      C@      K@     �z@     �S@     l�@     �k@     h�@     �u@      C@             �R@      e@      @      (@     �V@      @     `~@      G@     �r@      R@      @              B@     @U@      @      &@     �D@      @     �r@      <@     �^@      E@       @              2@      N@      �?      @      >@      @     `n@      4@     @U@      9@       @              .@      I@      �?      @      6@       @     �i@      4@     @S@      4@       @              @      $@                       @       @     �C@               @      @                      2@      9@       @      @      &@             �K@       @     �B@      1@                      ,@      6@              �?      @             �E@      @      7@      ,@                      @      @       @      @      @              (@       @      ,@      @                     �C@     �T@      @      �?      I@       @     �g@      2@     @f@      >@      @              A@      I@              �?      D@      �?     �S@      .@     �X@      8@      @              .@      ?@                      *@              C@      @      Q@      $@      @              3@      3@              �?      ;@      �?      D@      "@      >@      ,@                      @     �@@      @              $@      �?     �[@      @      T@      @       @              @      3@                      @             �R@              I@      �?       @              �?      ,@      @              @      �?     �A@      @      >@      @              (@      m@     x@      @@      E@     0u@     @R@     ��@     �e@     ~@     Pq@      ?@      (@     �d@     `m@      6@      ;@     �n@     �L@     �j@      b@     �h@     �h@      :@             �L@     @Q@       @      @     @S@      8@     @T@      G@      C@     �N@      "@              F@     �N@       @      @     �Q@      1@     �R@      >@      C@      I@      @              *@       @                      @      @      @      0@              &@       @      (@      [@     �d@      4@      7@      e@     �@@     �`@     �X@     �c@      a@      1@       @     �Z@     @d@      4@      7@      d@      <@     �`@     �W@     @c@     �`@      .@      @       @      @                       @      @      �?      @      @       @       @             �P@     �b@      $@      .@     �W@      0@     �u@      ?@     �q@      T@      @              D@     �Z@      �?      @     �M@      @     �q@      1@     `h@      L@      @             �A@     �Y@      �?      @      F@      @     �q@      0@     @g@     �J@      @              @      @                      .@               @      �?      "@      @                      ;@     �E@      "@      $@     �A@      "@     �P@      ,@     �V@      8@      �?               @      @               @      �?       @      $@      @      2@      "@                      3@     �B@      "@       @      A@      @     �L@      @      R@      .@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�3uJ�e@�	           ��@       	                    �?{ ���@�           L�@                          �<@I�;���@�           ��@                           �?�J86"Y@�           ��@������������������������       ��[(81�@           �z@������������������������       �_�F��@l            �e@                           �?�a`��@)            �L@������������������������       �bE��r @             2@������������������������       �V�HPx�@            �C@
                           @��cPx	@�           T�@                           �?�K�'N	@S           ��@������������������������       ��ɾ�͹	@i           ��@������������������������       ������a@�            0v@                          �9@�1�d�m	@�            �k@������������������������       �OX�]��@[             b@������������������������       �^{�ې�@*             S@                            �?�鄪�@3           ��@                           @�[��	�@@           ��@                          �6@�%,5�@�           ��@������������������������       �ռ�
@&           0}@������������������������       �ۘ�@h            �d@                           �?{��|�@�            �q@������������������������       ��R�rC[@S            �^@������������������������       �˖���@_             d@                           @��G�@�           ��@                           �?�"�=�@X           ��@������������������������       �����"�@�            �p@������������������������       ����;� @�            Pr@                            @�:ʱf@�            �k@������������������������       �oO:�:@J            �Z@������������������������       ��ĕ��@Q             ]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     0�@      ;@      Q@     �{@     �W@     ��@     `o@     x�@      u@      :@      *@     @k@      t@      7@     �H@     0t@     �Q@     �w@     @i@     �v@      m@      8@       @      S@      W@       @      "@     �R@       @     �c@      A@     `b@      J@      @       @      Q@     �S@       @      @      R@       @     �c@      <@     �a@      B@       @       @      L@     @P@       @      @     �J@      @     �W@      7@     �W@      ;@       @              (@      ,@               @      3@      @      O@      @      G@      "@                       @      *@               @       @               @      @      @      0@      �?              @      @                                      �?              �?      @                       @      @               @       @              �?      @      @      (@      �?      &@     �a@     �l@      5@      D@      o@     �O@     �k@      e@     �j@     �f@      5@      @     �^@     `h@      5@     �B@      j@     �H@     �g@      a@     �h@      d@      (@      @      Y@      b@      4@      @@      c@      D@     @\@     @X@     �b@     �\@      (@              6@      I@      �?      @      L@      "@      S@     �C@      I@     �G@              @      4@     �@@              @      D@      ,@      ?@      @@      0@      3@      "@      �?      0@      9@              @      ?@      $@      5@      (@       @      "@      "@      @      @       @                      "@      @      $@      4@       @      $@                     �T@     �l@      @      3@      _@      8@     ��@     �H@     `z@      Z@       @             �G@     �\@               @     �P@      *@     `t@      :@     �n@     @Q@                      :@     �T@              �?     �C@      "@      p@      0@     �c@     �E@                      1@     �M@                      ;@      "@     @j@       @      [@      =@                      "@      7@              �?      (@              G@       @     �I@      ,@                      5@     �@@              @      <@      @     �Q@      $@     @U@      :@                       @      (@              @      2@      @      :@      �?      D@       @                      *@      5@                      $@      �?      F@      "@     �F@      2@                      B@     �\@      @      &@     �L@      &@     �s@      7@     @f@     �A@       @              ;@     @T@              @      C@      @      n@      $@     @`@      7@                      6@     �F@              �?      2@       @     @X@      @      N@      1@                      @      B@              @      4@      @      b@      @     �Q@      @                      "@      A@      @      @      3@      @     �Q@      *@      H@      (@       @              @      4@       @      �?      *@      @      8@      @      8@      @       @               @      ,@       @      @      @       @     �G@      @      8@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Ϊ�A@�	           ��@       	                   �3@�?��@�           ��@                           �?5ɔ���@�           ��@                           @CH��&@�            r@������������������������       ��|."v�@�             m@������������������������       �j�"��@%             L@                           �?��m�Gf@           P{@������������������������       ��`��J@�             r@������������������������       �g����@^            �b@
                           �?����O^	@�           (�@                          �:@�6��?�@�            �x@������������������������       �z�q&~�@�            0r@������������������������       ����{kJ@B            �Z@                           �?9]̆�	@�           ��@������������������������       ��'v"?@�            �r@������������������������       �`&�?>�	@           ��@                           @��7b��@8           ��@                          �2@�j�s�@�           ��@                           @3��G��?           Pz@������������������������       �vI���a�?�            �s@������������������������       ��?i? @G             Z@                          �=@��p��@�           @�@������������������������       ���x�1�@�           (�@������������������������       �*~�9�@            �A@                           �?���u0A@Q           �@                          �0@*{�g\0@�            �h@������������������������       �N
�- �?             0@������������������������       ��\��@|            �f@                           @R�.��r@�            Ps@������������������������       �

�(^@�            �r@������������������������       ��ڇ8�E@             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     H�@      =@     �K@     �{@     �U@     8�@      i@     ��@     �w@      ?@      1@     @k@     �u@      5@      E@     �r@     @P@     �z@      f@     0w@      p@      <@      @      D@      [@      @       @     @R@      "@     @i@      L@     �a@     �S@       @      @      "@      H@       @             �@@      @     @U@      8@     �E@     �B@               @      @     �C@       @              ?@      @     �R@      1@     �B@      4@              �?       @      "@                       @       @      $@      @      @      1@                      ?@      N@      �?       @      D@      @     @]@      @@      Y@      E@       @              :@     �C@      �?      @      A@       @     �N@      8@     �N@      @@       @              @      5@               @      @       @      L@       @     �C@      $@              ,@     @f@     `n@      2@      A@     @l@      L@     @l@      ^@     �l@      f@      :@       @      >@     �R@      @       @     @R@       @     @S@      0@     �L@     �G@      �?              8@     �M@       @      @     �I@      @     �N@      $@      J@      5@      �?       @      @      0@      �?      �?      6@      @      0@      @      @      :@              (@     �b@      e@      .@      :@      c@      H@     �b@      Z@     `e@     @`@      9@             �@@     �C@       @      $@      C@      @      P@      1@     �K@      ?@      @      (@     �\@      `@      *@      0@     �\@     �E@     @U@     �U@      ]@     �X@      3@      �?     @Q@     @m@       @      *@     `b@      5@     �@      8@     @x@     �^@      @      �?     �F@     �c@       @      @     @T@       @     P}@      (@     Pq@     �R@      �?              "@     �M@      �?              .@              k@             �W@      ;@                       @     �D@      �?              "@             `e@             �P@      5@                      �?      2@                      @             �F@              <@      @              �?      B@     �X@      �?      @     �P@       @     �o@      (@     �f@      H@      �?      �?      @@      X@      �?      @      J@       @     �n@      (@      f@      G@      �?              @       @              �?      ,@              @              @       @                      8@     @S@      @       @     �P@      *@     �a@      (@     �[@      H@       @              @      B@               @      0@      @      S@      @     �G@      $@      �?                      @                      @               @                      @                      @      >@               @      *@      @     �R@      @     �G@      @      �?              3@     �D@      @      @      I@      $@     @P@      "@      P@      C@      �?              1@      D@      @      @      H@      @     @P@      "@     �O@      C@      �?               @      �?              �?       @      @                      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJz�%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?� ֥c@�	           ��@       	                   �;@�6Ӟ!|	@           ��@                           �?\xp�V!	@\           ��@                           �?S
�ܝ@B           �~@������������������������       �P����@@a            `b@������������������������       �z� ��;@�            `u@                           �?K5�	@           �@������������������������       ����?�@�            �p@������������������������       �����
@t           Ё@
                            �?�xU)�	@�            q@                           �?�O}��@.             R@������������������������       ��]��G#@             8@������������������������       �����@             H@                            �?σk �
@{             i@������������������������       �܈�Y�@)            �M@������������������������       �%N���	@R            �a@                           @�>K�XQ@�           �@                           �?Ȫ�o@h           �@                            �?&rʩA�@s            �g@������������������������       ���y4@%            �N@������������������������       ��,U�@N            �_@                            @z���@�            Pv@������������������������       ��
r8��@�            �o@������������������������       ��*vO7�@N            @Z@                           �?_=���t@;           ��@                           @�aR��� @j           ��@������������������������       ����
�?�            �x@������������������������       ��?�w�@~            `i@                          �7@�Lۻ�p@�           X�@������������������������       ��� �b@"           Ћ@������������������������       �ߦ�x`@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �q@     �@      B@     �G@     pz@     @Q@     ��@     �j@     Ȉ@     @w@      :@      6@     �d@     �l@      <@      C@      k@      G@     �n@     @`@     `o@     @i@      5@      (@      a@     �g@      7@      =@     �f@      =@      l@     @[@     �l@     �a@      4@      �?      A@     �R@       @      ,@     �Q@      @     @Z@     �C@      U@      M@      @              (@      2@                      5@              D@      @      E@      "@      �?      �?      6@      L@       @      ,@      I@      @     @P@     �A@      E@     �H@      @      &@     �Y@     �\@      5@      .@      \@      :@      ^@     �Q@      b@     �T@      0@             �A@     �D@      @      @      :@      �?     �M@      1@      J@      3@      @      &@      Q@     @R@      .@      $@     �U@      9@     �N@     �J@      W@      P@      (@      $@      <@     �E@      @      "@      A@      1@      5@      5@      7@     �N@      �?              @      .@                      &@      �?      @       @      @      4@      �?                      @                       @      �?      @      @      @      �?                      @       @                      "@              @      @      �?      3@      �?      $@      9@      <@      @      "@      7@      0@      ,@      *@      1@     �D@              @      $@      @       @      @      @       @      @       @      @      1@              @      .@      7@      @      @      4@      ,@      &@      @      ,@      8@                      ^@     �s@       @      "@     �i@      7@     �@     @U@     ��@     @e@      @              C@     �T@       @      @      M@       @     `b@     �D@     �Z@      L@       @              3@      .@              �?      0@             �Q@      @      G@      ,@       @               @      @              �?      @              5@              7@      @       @              1@      &@                      (@             �H@      @      7@      $@                      3@      Q@       @       @      E@       @     @S@      B@     �N@      E@                      (@     �C@       @      �?     �C@      @     �L@      4@     �H@      :@                      @      =@              �?      @      �?      4@      0@      (@      0@                     �T@     �l@      @      @     �b@      .@     x�@      F@     0{@     �\@      @              4@     �R@      �?      �?      9@      @     @s@      $@     �_@      8@      �?              *@      E@                      $@      @     @m@       @      S@      (@                      @      @@      �?      �?      .@      �?     �R@       @     �I@      (@      �?              O@     �c@      @      @     �^@      "@     �w@      A@     @s@     �V@       @             �C@     �_@      @      @      S@      @     �s@      (@     �n@     �M@       @              7@      ?@      �?       @     �G@       @     �N@      6@      P@      ?@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?w�mw@�	           ��@       	                    �?�g�(N\	@           ؙ@                          �<@Pٚ�C@1           �~@                           �?p�R��`@           p{@������������������������       �F�ɛ��@�            �i@������������������������       �c@��mV@�            `m@                           �?.�À@!             K@������������������������       ��7����@             2@������������������������       ��:��0@             B@
                          �<@OlI3��	@�           $�@                           �?�g:��	@�           ��@������������������������       ��_DX��@�            �w@������������������������       �	����O
@�           ��@                           @U&���	@_             b@������������������������       �*�%WQ@             @@������������������������       �d�a�6@H            @\@                          �5@� �dm+@�           ��@                           @SǻGu_@w           ��@                            �?As� ��@d           ��@������������������������       ����@�            �t@������������������������       ����&l@�            �l@                           @�����@           ��@������������������������       �r�qhq�@�           ��@������������������������       �Ĭ���@$             L@                          �<@�?�	�/@,           ��@                          �9@ٖ1c�@�           0�@������������������������       ��W���$@W           X�@������������������������       ��Z�g�Y@|            `g@                           @���V@Y            `a@������������������������       ���`�w	@             D@������������������������       �^b�g>�@=            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `r@     ��@     �C@     �O@     p}@     @T@     h�@      l@     �@     �u@      @@      1@     �d@      m@      @@      E@     �p@      E@     �m@      a@     Pq@     �f@      8@              I@      N@              @     @S@      @     �Z@      ?@     @[@     �B@       @             �E@      M@               @     �P@      @     @Z@      ;@     �Y@      4@       @              4@      2@                      C@      @      H@      .@     �D@      ,@      @              7@      D@               @      =@             �L@      (@     �N@      @      @              @       @              @      $@               @      @      @      1@                      @      �?                       @               @               @      @                       @      �?              @       @                      @      @      &@              1@     �\@     �e@      @@     �A@      h@     �A@     @`@     @Z@      e@      b@      0@      ,@     �Y@      c@      ?@      <@     `e@      7@     @^@     �V@     @c@     �\@      ,@      �?     �@@      Q@      @       @     @Q@      @      P@      :@     �J@     �G@       @      *@     �Q@      U@      <@      4@     �Y@      1@     �L@      P@     @Y@      Q@      (@      @      &@      4@      �?      @      5@      (@      "@      .@      ,@      >@       @       @       @       @      �?      @      @      @      �?       @      @      @       @      �?      "@      2@              @      2@      "@       @      *@      "@      9@              @     @`@     �r@      @      5@     @i@     �C@      �@     @V@     h�@     �d@       @             @P@      g@      @       @     @V@      .@     `�@      D@      u@     �R@      @              B@      V@      �?      �?     �A@      *@     @h@      ;@      `@      C@      �?              6@      J@              �?      1@      $@     @`@      0@     @R@      *@                      ,@      B@      �?              2@      @      P@      &@     �K@      9@      �?              =@     @X@      @      @      K@       @     �v@      *@      j@     �B@      @              :@     �W@      @      @     �I@       @     �u@      *@     `h@      8@      �?              @      @              �?      @              2@              *@      *@       @      @     @P@      ]@       @      *@     @\@      8@     �j@     �H@     �g@     �V@      @      @     �G@      Z@       @      $@     @T@      4@     `h@      E@      d@     �R@      @      @      B@     @S@      �?      "@     �P@      .@      b@      ;@     �Z@     �P@      @              &@      ;@      �?      �?      .@      @      I@      .@      K@       @                      2@      (@              @      @@      @      1@      @      <@      1@      �?              @      @               @      @      @       @      @      @       @      �?              *@      @              �?      ;@      �?      .@      �?      9@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJa"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�b�;@�	           ��@       	                    �?�c^k,�@v           ��@                          �6@[i9"P@�           ��@                          �4@�*u�,�@           �{@������������������������       ��t��@�            �t@������������������������       �MDpyz@@            @[@                            @h4��@�            �o@������������������������       ��F���N@k            @d@������������������������       �,�K�S�@=             W@
                           �?�����`	@�           �@                            @�����@I            �^@������������������������       �,�N�.�@)             O@������������������������       ���0�\V@             �N@                           �?cEE��0	@r           (�@������������������������       ��3��)�	@�           ��@������������������������       �1:}onV@�            `w@                           @��5 U�@6           8�@                          �4@�|N�S<@�           ��@                            @�z� @�           �@������������������������       �q�p^{ @�           p�@������������������������       �D�r�8��?4             U@                            @L����@0            ~@������������������������       ���H��@           �y@������������������������       ��o/���?+            @P@                           �?�	�M�@N           `�@                          �:@\{=�\@�            pq@������������������������       ��#�N�^@�             m@������������������������       ��NZY�@             G@                            �?�U���@�            Pq@������������������������       ������ @&            �O@������������������������       ��*�v�@�            �j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     pr@     ��@      ;@     �L@     @|@     @T@     h�@      k@     (�@     pv@      8@      .@     �k@      s@      6@     �F@     �s@     �N@     �w@      f@     @v@     �o@      2@      �?     �S@     @V@       @      $@      S@       @      h@     �D@     �a@     �L@      @              I@      I@              @     �E@       @     �b@      :@     �W@      7@                      <@      E@                      D@       @     @Z@      4@     @S@      1@                      6@       @              @      @              F@      @      1@      @              �?      =@     �C@       @      @     �@@             �E@      .@      H@      A@      @      �?      5@      ;@              @      1@              >@      @      ;@      :@      @               @      (@       @      @      0@              *@       @      5@       @              ,@     �a@      k@      4@     �A@     @n@     �M@     `g@      a@     �j@     �h@      .@       @      4@      ,@              (@      ,@      @      �?      ,@      2@      5@      �?              @       @              @       @       @              @      .@      ,@      �?       @      *@      (@              @      @      @      �?      @      @      @              (@     �^@     `i@      4@      7@     �l@     �J@     @g@     �^@     �h@     �e@      ,@      (@     �X@     �a@      1@      6@     �d@      B@     @[@      V@      a@     �a@      ,@              8@      O@      @      �?      O@      1@     @S@      A@      N@      A@                     �R@     @l@      @      (@     �`@      4@     ��@     �C@     |@     �Z@      @              H@     �a@       @      @     �T@      $@     p@      0@     �s@      O@      @              :@     �S@               @      @@       @     �u@      @      h@      7@                      6@      R@               @      >@       @     �s@      @     �b@      6@                      @      @                       @              :@      �?     �E@      �?                      6@      P@       @      �?     �I@       @     �c@      $@     @^@     �C@      @              4@      P@       @      �?     �H@      @     @_@      $@      Y@     �A@       @               @                               @      �?      A@              5@      @      �?              :@     �T@      @      "@     �I@      $@      e@      7@      a@      F@      @              "@      A@       @      "@      :@      @     �W@      "@     @Q@      7@                      @      >@       @      "@      8@       @     @S@      @     �N@      5@                      @      @                       @       @      1@      @       @       @                      1@     �H@      �?              9@      @     �R@      ,@     �P@      5@      @              @      @                      @      @     �A@      @       @                              ,@      F@      �?              3@      @     �C@      &@     �M@      5@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?>��"@�	           ��@       	                     @y��n|@           ��@                          �8@)���?�@F           ��@                          �2@t)��[u@�           x�@������������������������       �T���� @�             s@������������������������       �5���@           �{@                          �<@�y��i@q             f@������������������������       �{}|�4@@            �Y@������������������������       �����6@1            @R@
                           �?td�v�@�            �t@                          �9@�X`�"@f            �c@������������������������       ��<o��@N            @^@������������������������       ��Jv@             B@                          �:@(�s��@l            �e@������������������������       �kc��O @a            �c@������������������������       ���	M�1@             0@                           @��AI$@�           ��@                          �5@P8�~�@^           0�@                            @��#�@c           Е@������������������������       �e�Ƃ�@w           ��@������������������������       ���Y�s@�            �w@                           @��]��@�           ��@������������������������       �\�=k�k	@�           �@������������������������       ��HZ�H@           pz@                            �?
�IG��@.            �Q@������������������������       �]�d�@             4@                          �4@��=��@#            �I@������������������������       �Nɱ���@
             ,@������������������������       �j�v%�@            �B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     p@     ��@      =@     �M@     0|@     @Q@     ��@      l@     8�@      x@      >@             �Q@      f@      �?      @     �W@      &@      |@      H@     t@     @S@      @             �G@      `@      �?       @     �P@      $@     u@      :@      p@     �G@      @             �B@     �Y@      �?       @     �G@      @     �r@      (@     �i@      >@      @              *@      @@              �?      1@             @c@      @     �P@      0@       @              8@     �Q@      �?      �?      >@      @     �b@       @     �a@      ,@      �?              $@      :@                      3@      @      A@      ,@     �H@      1@      @              @      ,@                      &@      @      9@       @      @@       @       @              @      (@                       @              "@      @      1@      .@       @              7@      H@               @      =@      �?     �[@      6@     @P@      >@                      "@      2@               @      8@      �?     �J@      "@      <@      *@                      "@      .@                      &@      �?      F@       @      5@      (@                              @               @      *@              "@      �?      @      �?                      ,@      >@                      @              M@      *@     �B@      1@                      (@      =@                      @              L@       @     �B@      *@                       @      �?                       @               @      @              @              1@     `g@     �v@      <@     �K@     @v@      M@     ��@      f@     0�@     0s@      7@      .@      f@     Pv@      ;@     �K@     `u@     �K@     ��@     @d@     �@     �r@      4@       @      J@      i@      &@      <@     @d@      5@     `w@      T@      t@      `@      "@      �?      D@     `b@       @      2@     �Z@      "@     Pr@     �L@      n@     �Y@      @      @      (@     �J@      "@      $@      L@      (@     @T@      7@     @T@      ;@      @      @     @_@     �c@      0@      ;@     �f@      A@     �g@     �T@     `g@     �e@      &@      @      W@     �[@      &@      2@     @`@      >@     �S@     �P@      U@     @_@      &@             �@@      G@      @      "@      I@      @     �[@      .@     �Y@      H@               @      $@      @      �?              ,@      @      @      ,@      "@      @      @              @      @      �?              �?                      @       @                       @      @      @                      *@      @      @       @      @      @      @      �?              @                       @               @              �?       @      @      �?      @      �?                      &@      @      �?       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>�W"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @ڰ�*�@�	           ��@       	                   �8@���
		@�           ��@                           �?h(�B2@�           @�@                           �?|� w_@.           �}@������������������������       �����@�            @j@������������������������       �~AJ�@�            �p@                           @5��#�@�           Б@������������������������       ������@�           X�@������������������������       �����@             >@
                          �:@Lso��
@�           �@                           @�'�	@�            @k@������������������������       ��U)D �@i            �d@������������������������       �Bɾޅ�@%             K@                          �<@ �Io�	@           �z@������������������������       �˚�`J	@_            @d@������������������������       �:m˚>%	@�            `p@                            @d'�Fz�@           ܙ@                           �?�:S�@s           ��@                           @긲t@"           �|@������������������������       ��'�q��?�            �s@������������������������       ���/<�@[            �a@                           @��Dg@Q           �@������������������������       �5��&�@           ��@������������������������       ���J@E            �[@                           �?R̞Y�C@�            �p@                           �?t�K�k�?;            �U@������������������������       �w����Q�?!             F@������������������������       �n�A����?             E@                           @�࿎@p             g@������������������������       ��D��/@@            �Y@������������������������       ��K8ܥ%@0            @T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     @s@     �@     �A@     �I@     @|@      V@     ��@     `k@     ȇ@     �w@      B@      4@     �l@     �u@      8@      E@     �t@     �Q@     �u@     @f@     �v@     �p@      >@      @     �c@     `o@      ,@      ;@     �n@      C@     r@     �]@     s@      c@      .@              B@     �P@      @       @      M@      �?     `a@      6@     �[@     �@@                      0@      ;@      @              B@      �?      P@      *@      @@      ,@                      4@      D@               @      6@             �R@      "@     �S@      3@              @      ^@      g@      @      9@     �g@     �B@     �b@      X@     @h@     �]@      .@      @     �\@     �f@      @      9@     `f@      B@     �b@     �W@      h@      ]@      $@       @      @       @                      "@      �?      �?      �?      �?      @      @      .@     @R@     �X@      $@      .@      U@      @@      O@      N@     �N@     @]@      .@              >@     �G@      @      @      ;@      $@      3@      5@      3@      8@      &@              :@      @@              @      3@      "@      ,@      .@      0@      7@      @              @      .@      @       @       @      �?      @      @      @      �?      @      .@     �E@     �I@      @       @     �L@      6@     �E@     �C@      E@     @W@      @      (@      *@      1@      @              5@      @      8@      *@      :@      <@      �?      @      >@      A@      @       @      B@      2@      3@      :@      0@     @P@      @      @     �S@      l@      &@      "@     �^@      2@     �@     �D@     �x@     �[@      @      @     �P@     �i@      @      @     @Y@      ,@     ��@      C@     �s@     @W@      @              (@     @Q@      �?              8@      @      l@      @      X@      1@       @              &@      D@                      (@       @     @f@      @      N@      "@                      �?      =@      �?              (@       @      G@      @      B@       @       @      @      K@      a@      @      @     @S@      $@      s@      ?@     �k@      S@      @      @     �C@      `@      @      @     �Q@      @     �p@      <@     �i@     �O@      �?              .@      "@       @      �?      @      @     �D@      @      .@      *@       @              *@      2@      @       @      5@      @     �Z@      @     �S@      1@      �?              @      @                      �?             �K@              8@                              @       @                                      ?@               @                                      �?                      �?              8@              0@                              $@      .@      @       @      4@      @      J@      @     �K@      1@      �?              @       @                      *@      �?      A@              D@      @      �?              @      @      @       @      @      @      2@      @      .@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJH��7hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?5��ˁJ@�	           ��@       	                    �?�K:�@�@�           �@                           @��T��'@�            �u@                          �;@L]!m�@y            �i@������������������������       �����@n             h@������������������������       ��悛@             ,@                          �4@�����?Y            �a@������������������������       �&a�mg2�?9             X@������������������������       ��L��K|@             �F@
                           @��!@^�@�           8�@                          �4@@�X��,	@            z@������������������������       �E�o�@c             c@������������������������       ��'�P�	@�            �p@                           @5{J;C�@�            Pp@������������������������       �,i�#`�@8            @U@������������������������       ��U�X��@u             f@                           �?�X!�f@           ��@                           �?r�0ƚ@           X�@                            @I��@           p}@������������������������       �7}?\�@�            pq@������������������������       �0���!~@l             h@                            �?K��A��@�            @w@������������������������       �M�Nô)@b             b@������������������������       � y���@�            �l@                           @P���)6@�           �@                           �?��ԕ	z	@�           ��@������������������������       ��O��J�	@�            �x@������������������������       ��@
�� 	@�           ��@                           @���5/@;           Ȍ@������������������������       �&ށ���@�           ؃@������������������������       �b}���=@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@     �@@     �M@      |@     @S@     ��@     �k@     H�@     �u@      :@      �?     @T@     �_@      @      $@     @\@      9@     �r@     �S@     @i@     @S@       @      �?      3@     �E@      �?              :@      @     �a@      &@     �U@      .@      �?      �?      3@      >@                      0@       @      J@      &@      P@      &@      �?              1@      ;@                      .@      �?      J@      &@     �O@      @              �?       @      @                      �?      �?                      �?      @      �?                      *@      �?              $@      �?     @V@              7@      @                               @                                     @Q@              1@       @                              @      �?              $@      �?      4@              @       @                      O@      U@      @      $@     �U@      6@      d@     �P@     �\@      O@      @             �D@      J@      @      $@      P@      5@      O@     �L@     �L@      F@      @              (@      .@                      7@      @     �C@      3@      9@      ,@       @              =@     �B@      @      $@     �D@      2@      7@      C@      @@      >@      @              5@      @@                      7@      �?     �X@      $@      M@      2@                      (@      .@                      @              :@      @      ,@      $@                      "@      1@                      2@      �?      R@      @      F@       @              3@     @k@      {@      =@     �H@     u@      J@     (�@      b@     ��@     �p@      2@              Q@     @]@       @      &@      T@      @     �q@      6@     �h@     �K@       @              F@     @P@       @      "@     �I@             �c@      0@     �W@      >@      �?              :@     �D@      �?      @      ?@             �Y@      $@      I@      *@      �?              2@      8@      �?      @      4@              L@      @     �F@      1@                      8@      J@               @      =@      @      `@      @     @Y@      9@      �?              @      3@                      @      @     �G@      �?      I@      ,@                      2@     �@@               @      9@             �T@      @     �I@      &@      �?      3@     �b@     �s@      ;@      C@     p@     �H@     `z@     �^@     �y@     �j@      0@      1@     �Y@     �f@      .@      ;@     �e@     �E@     �a@     @Z@      e@     `a@      &@      "@     �D@     @Q@       @      "@     �J@      2@      I@     �B@      G@     �J@      @       @     �N@     �[@      @      2@     �]@      9@      W@      Q@     �^@     �U@      @       @      H@      a@      (@      &@     @U@      @     �q@      2@     @n@     �R@      @       @      =@     �X@       @      @     �J@      @      l@      "@      e@      C@      @              3@     �C@      $@      @      @@      @      L@      "@     @R@     �B@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ%D�fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�Bx                             �?!�Pc]@�	           ��@       	                     �?�?���1@�           �@                          �8@	���5@�            �t@                           �?0W�ڇl�?�            �p@������������������������       �����@5            �V@������������������������       ���l�Z��?l            @f@                           �?#��K�@*            �P@������������������������       ���< �@             >@������������������������       ����p7�@             B@
                          �<@/�+���@'           h�@                           �?�װ��@�           ��@������������������������       �
��3�@�            �q@������������������������       �͊a��@D           0�@                            �?y��!<[@3            �S@������������������������       �z�s����?             B@������������������������       �X)�-��@             E@                           !@9�[X@�           �@                           �?�p���B@�           �@                          �7@<�*���	@~            �i@������������������������       �ٵR�]@Q            �`@������������������������       ����@-            @Q@                           @�g�_ @           T�@������������������������       �qQ��YV	@�           p�@������������������������       ����2��@�           8�@������������������������       �I��y�}@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B`	        ?@     �p@     P�@      ?@     �K@     �y@      X@     �@     @k@     h�@     @w@      <@      @     �S@      d@      �?      *@     �V@      @     �|@     �E@     0q@      U@      @      @      &@     �F@              �?      @@      �?     �b@      @     �Q@      .@                      @      A@              �?      7@             �`@       @     �O@      @                      @      (@                      &@              <@       @      ?@      @                              6@              �?      (@             �Z@              @@      @              @       @      &@                      "@      �?      0@       @       @       @              @      @      @                       @              @       @       @      @                      @      @                      @      �?      $@              @       @                     �P@     �\@      �?      (@     �M@       @     s@     �C@     �i@     @Q@      @             �M@     �Z@      �?       @     �I@       @     �r@      A@     �g@      G@      @              9@     �E@      �?      @      8@       @     �P@      4@      P@      <@      @              A@      P@              @      ;@             �l@      ,@     �_@      2@      �?               @       @              @       @              "@      @      *@      7@                      @                       @                      @       @      @      4@                      @       @               @       @              @      @       @      @              <@      h@     �x@      >@      E@      t@     @W@     ��@     �e@     Ѐ@      r@      8@      <@     �g@     �x@      >@      E@     �s@     �T@     ��@     �e@     ��@      r@      6@      @      *@      8@              ,@      ;@      (@      6@      3@     �E@      5@      @       @      @      5@              "@      ,@      &@      6@      @      =@      0@              @      @      @              @      *@      �?              ,@      ,@      @      @      6@      f@     w@      >@      <@     @r@     �Q@     H�@     �c@     �~@     �p@      3@      6@     ``@     �j@      5@      4@      g@     �J@     �j@     �`@      n@     �f@      2@              G@     `c@      "@       @     �Z@      1@      u@      5@     @o@     �U@      �?              @      �?                      @      &@                      @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{�`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Q�.�a@�	           ��@       	                   �6@���h�L@(           ��@                          �1@/':�Sv@           @�@                          �0@�m�PN* @�            �n@������������������������       ��)�,�?6            @T@������������������������       ���p|[l @o            �d@                          �3@��Q@w           ��@������������������������       ��Sq",@�            `s@������������������������       �Ғ1_�@�            �q@
                            @�4^��@            z@                           �?(7T-��@�            s@������������������������       �$�çS@[            �a@������������������������       ����̔@i            �d@                          �7@E��:@H            �[@������������������������       ���(r�T�?             1@������������������������       ����^�@;            �W@                          �7@�}�1D
@}           ¤@                            @�{�@�@e           �@                          �4@!�\���@:           \�@������������������������       �&�R^Z@           ȉ@������������������������       ���=�&�@(           �}@                           @�6'�y�@+            @������������������������       �G6�F@�            `v@������������������������       �1>���i@O            @a@                           �?|[�C�k	@           Њ@                            �?`���	@           �}@������������������������       �����.�@�             l@������������������������       �C�)5�	@�             o@                           �?�K���K@�            x@������������������������       ����5C�@l            `f@������������������������       �d/zM@�            �i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     ��@      ;@      E@     �x@     @P@     ,�@     @o@     @�@     pw@     �@@      �?     �V@     `d@      @      @      V@      @     0}@     �J@      r@     @T@      @             �I@      \@              @      E@      �?      w@      :@     �g@     �E@      @              $@      8@              �?      @             �^@      @     �P@       @      @                      @                      @             �E@       @      6@      @                      $@      1@              �?      @              T@      �?     �F@      @      @             �D@      V@              @     �A@      �?     �n@      7@     �^@     �A@                      7@      E@              �?      ,@              ]@      (@     �S@      8@                      2@      G@               @      5@      �?      `@      &@     �F@      &@              �?      D@     �I@      @       @      G@      @     �X@      ;@      Y@      C@      @      �?      >@     �E@      @             �@@      @      N@      0@     �S@      A@      @      �?      1@      4@                      *@      �?      @@      "@      ;@      4@                      *@      7@      @              4@      @      <@      @     �I@      ,@      @              $@       @       @       @      *@             �C@      &@      6@      @                                                       @              @               @      �?                      $@       @       @       @      &@             �@@      &@      ,@      @              1@     @j@     y@      6@      B@     0s@      N@     ��@     �h@     0�@     `r@      ;@      @      b@     �q@      (@      7@      g@      9@     �|@     @V@     �x@     `e@      *@      @     �X@      h@       @      3@      a@      .@      v@     �P@      r@     �\@       @      �?      J@      [@      @      @      Q@      @     �p@      F@     `h@     �R@      @       @      G@      U@      �?      0@      Q@      &@     �V@      6@     �W@      D@      @      @     �G@     @V@      @      @     �H@      $@     �Y@      7@     �Y@     �L@      @      @      B@     �Q@      @      @     �E@      $@     �L@      6@      O@     �F@      @              &@      3@      �?              @             �F@      �?     �D@      (@       @      &@     @P@      ^@      $@      *@     �^@     �A@      \@      [@     @_@     �^@      ,@      "@      D@      M@       @       @      N@      ;@      E@     �S@      E@     �U@      ,@      @      .@      :@       @      @      3@      4@      0@     �K@      4@      D@      @      @      9@      @@      @      @     �D@      @      :@      7@      6@     �G@       @       @      9@      O@       @      @      O@       @     �Q@      >@     �T@      B@               @      "@     �@@              @      >@       @      9@      $@      E@      6@                      0@      =@       @      �?      @@      @     �F@      4@     �D@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��9ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@7��'@�	           ��@       	                    �?s]��Á@p           ̛@                           �? �+m�U@�           ��@                           �?�/�@y            �f@������������������������       �{��N�@3            �S@������������������������       �>м�E�@F             Z@                           �?������?#           �}@������������������������       ��47
`n�?�             o@������������������������       ����j�?�             l@
                           @ԫR���@�           ��@                           �?��E^b�@g           X�@������������������������       �����o@�            @w@������������������������       �F��0.@v            �f@                           �?�PTNT�@m           ��@������������������������       ���iD�3@�            �r@������������������������       ��:ǅ�@�             q@                           �?���>f@O           ��@                          �<@%uMv��@z           p�@                            �?���r��@>           `~@������������������������       �����@U            �^@������������������������       �E�z԰@@�            �v@                            @���ɨ�@<             Z@������������������������       �J�O(<R@*            �R@������������������������       �����@             =@                           @ ���	@�            �@                          �9@7W<�:	@h           ��@������������������������       ���YvQ@�           0�@������������������������       �����
@�            �t@                          �:@"K�)�@m           ��@������������������������       ��r��@�            `y@������������������������       �$�z�L4@n            �c@�t�b��     h�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     �@      6@     �F@      {@      W@     ��@     `j@     ��@      v@      >@       @     @Z@     �l@      @      ,@     �d@      .@     X�@      N@     �v@      _@       @              6@     �R@              @      C@       @      u@      1@     �_@      ?@      @              @      >@              �?      2@       @     �P@      *@      ?@      .@                      �?      ,@                      @              ?@      @      4@      @                      @      0@              �?      *@       @     �A@      "@      &@      &@                      .@      F@              @      4@              q@      @     �W@      0@      @              @      6@              @      .@             �a@      @      F@      *@                      &@      6@                      @              `@             �I@      @      @       @     �T@     �c@      @      "@     �_@      *@     �u@     �E@      n@     @W@      @       @     �G@      T@      @      @     �W@      $@     �[@     �B@     �X@      O@      @       @     �C@     �C@      @      @     @Q@       @     �N@      :@     @Q@      F@      @               @     �D@                      9@       @     �H@      &@      =@      2@                      B@     @S@       @      @      @@      @     `m@      @     �a@      ?@                      4@      ?@       @      @      6@      �?      ^@      @     �R@      2@                      0@      G@                      $@       @     �\@       @      Q@      *@              &@     �h@     �s@      .@      ?@     �p@     @S@     �x@     �b@     0z@     �l@      6@              J@      W@      �?      @     �L@      (@      e@      8@      `@     �H@                     �F@     �S@      �?      @      F@      (@     @c@      .@      ]@      2@                      &@      2@      �?       @      ,@      @     �A@      �?      <@      @                      A@      N@              �?      >@      @     �]@      ,@      V@      (@                      @      ,@               @      *@              .@      "@      *@      ?@                      @       @                      @              &@      @      $@      <@                      �?      @               @       @              @       @      @      @              &@      b@     �k@      ,@      :@     �j@     @P@     �l@     �_@      r@     �f@      6@      &@     �X@      ^@      "@      3@     `a@      K@      b@     �M@     �h@     �[@      1@      @     �O@     �S@      @      ,@     @W@      8@     �]@      9@     @a@     �R@      "@      @      B@     �D@      @      @      G@      >@      :@      A@     �N@     �A@       @              G@     �Y@      @      @     �R@      &@      U@      Q@     �V@     �Q@      @              ?@     �V@      @      @     �I@      @      M@      I@     �Q@      A@      @              .@      &@              @      7@      @      :@      2@      5@     �B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�)$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�O:4@�	           ��@       	                     @w�ɝS�@�           t�@                           @X��\�@�           ��@                           @�f5V#.@           �y@������������������������       ��˜~��@�             t@������������������������       ��U�W�@=            �V@                           @��xy.@�           �@������������������������       �k�֢� @/           �~@������������������������       ��F��@U            @^@
                           �?�����@�            �y@                           @)|�-Ⱥ@]            �c@������������������������       ��5w���@C            �\@������������������������       �ΟH�b��?             F@                           @�0s��@�             p@������������������������       �̨�f��@r             g@������������������������       �[~��Q@@*             R@                          �9@��-5@'           X�@                           �?:�rΆ@E           �@                           �?��v�`�@:            }@������������������������       �RGZ�@�            Pp@������������������������       ��%&�l9@�            `i@                            @����0@           Г@������������������������       ��)k� �@5           P�@������������������������       ��\Ne�J@�            �v@                          �;@���h'	@�           @�@                          �:@�hs�,@�            s@������������������������       ���+~@f            �d@������������������������       ��"��@]            @a@                           �?z ��m	@           p{@������������������������       ���k�@J            �[@������������������������       ����ۗ�	@�            �t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     ��@      ?@     �G@      ~@     �R@     ��@     �h@      �@     �u@      =@      @     �U@     �g@      @      (@     ``@      &@     �~@     �H@     0v@      Y@       @      �?      I@     �`@      @      @     @T@      @     w@      >@     �p@      R@       @      �?      <@     �J@      @      �?      I@      @      V@      :@     �\@      E@      �?              :@      @@       @      �?      B@      @     �P@      2@     @X@     �B@              �?       @      5@      �?              ,@              5@       @      1@      @      �?              6@     �T@      @      @      ?@             �q@      @     @c@      >@      �?              4@     �P@      �?              4@              n@      @     �]@      3@                       @      .@       @      @      &@              D@      �?     �A@      &@      �?      @      B@      L@      �?       @      I@      @     �]@      3@     �U@      <@                      1@      ,@              @      $@      �?      Q@      @      C@      @                      1@      *@              @      $@      �?     �B@      @      :@      @                              �?                                      ?@              (@                      @      3@      E@      �?      @      D@      @     �I@      0@     �H@      7@               @      $@      ;@      �?       @      =@      �?     �B@      ,@     �E@      2@               @      "@      .@              @      &@      @      ,@       @      @      @              2@     �j@     pw@      8@     �A@     �u@      P@     �~@     �b@     �}@      o@      ;@      @      b@     @q@      1@      9@     p@      >@     0x@      U@     �u@      a@      4@             �D@      W@      @      @     �H@       @     @a@      (@     �Y@      3@      �?              5@     �E@       @      @      @@              W@      $@     �G@      $@                      4@     �H@      �?              1@       @      G@       @      L@      "@      �?      @      Z@      g@      ,@      5@      j@      <@      o@      R@     �n@     �]@      3@       @     @S@     �_@      @      5@      a@      5@      i@     �J@     �e@     �T@      $@      @      ;@     �L@      $@              R@      @     �H@      3@      R@     �A@      "@      &@     �Q@     �X@      @      $@      W@      A@      [@      P@     @`@      \@      @              9@      A@       @       @     �B@      0@     �I@     �@@     �P@      B@      @              .@      6@       @      �?      2@      .@      9@      .@      C@      ,@       @              $@      (@              �?      3@      �?      :@      2@      <@      6@      �?      &@     �F@     @P@      @       @     �K@      2@     �L@      ?@      P@      S@      @      �?      "@      .@              @      (@              :@      "@      3@      1@              $@      B@      I@      @      @     �E@      2@      ?@      6@     �F@     �M@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��9OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@Q���*@�	           ��@       	                    @`8��j@�           �@                           @�jF�@>           �@                          �1@���w�@�            y@������������������������       �����ʉ@�            `k@������������������������       ��^�7�@m            �f@                           @�X�i2:@K             [@������������������������       �(T��]�@9            �T@������������������������       ���� �@             :@
                           @��<Ƭ @c            �@                           @�%���?�            0t@������������������������       �ms��T�?6            �U@������������������������       ��A�}���?�            �m@                            �?v�S���@�            p@������������������������       �|=&�?              J@������������������������       ��x*���@�            �i@                          �<@�R�\@+           �@                           �?`=yR��@W           t�@                            @�/�\�@�           �@������������������������       ��:���L@>           �}@������������������������       �;�j}n@�            �h@                            �?�,fn�@�           \�@������������������������       ��k�S�@I           �@������������������������       �Z�s�w@K           t�@                          @A@t�u�J@�            �t@                           �?��%p��@�             s@������������������������       �(Gi�ε@<            @W@������������������������       ��Bal�@�            `j@                           @��<rD�@             >@������������������������       �JE}�u) @             ,@������������������������       �|R��>@             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �p@     H�@      4@      H@     �{@     @U@      �@     �l@     h�@     w@      @@       @      F@     �a@              @     �Y@      @     p|@      F@     �j@     �S@       @       @      >@      P@              @     �R@       @     �b@      B@     @W@      K@      �?              5@      C@               @     �O@      �?     @_@      7@     �T@      G@                      @      7@              �?      9@             @T@      (@      J@      2@                      ,@      .@              �?      C@      �?      F@      &@      >@      <@               @      "@      :@              �?      (@      �?      8@      *@      &@       @      �?       @      @      6@              �?      @              5@      (@      @      @                      @      @                      @      �?      @      �?      @      @      �?              ,@      S@              �?      ;@       @      s@       @     @^@      8@      �?              @     �C@                      @       @     �i@      @      H@      "@      �?               @      3@                               @      I@              (@       @                      @      4@                      @             `c@      @      B@      @      �?              @     �B@              �?      4@             @Y@      @     @R@      .@                      �?      @              �?      @              >@               @      @                      @      A@                      .@             �Q@      @     @P@      &@              2@     �k@     �{@      4@      F@     Pu@     @T@     �@     `g@     ��@     0r@      >@      ,@     �h@     px@      0@      B@     �r@     �Q@     (�@     @c@     @�@     �j@      >@             �F@     �Y@       @      @     �M@      @      j@      =@     @f@     �C@      @              ;@     @Q@                      C@      @      c@      5@     ``@      ;@      @              2@     �@@       @      @      5@             �K@       @     �G@      (@              ,@      c@     r@      ,@     �@@      n@      P@     Pu@     @_@     `u@     �e@      ;@       @      J@     �R@       @      &@     �L@      2@     @V@     �J@     �U@     �K@      @      (@      Y@     �j@      (@      6@      g@      G@     �o@      R@     �o@     �]@      5@      @      :@      K@      @       @     �D@      $@      <@     �@@     �G@     �S@              @      6@     �H@               @     �C@      @      <@     �@@      E@      R@                       @      *@              @      "@              &@      0@      *@      :@              @      4@      B@              @      >@      @      1@      1@      =@      G@                      @      @      @               @      @                      @      @                      �?      @                      �?                              @      @                      @       @      @              �?      @                       @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ92hyhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?B�yA1 @�	           ��@       	                    �?<�r�Ú@           h�@                           �?��"W�@-           p}@                          �3@��n ��@�            �j@������������������������       ����?��@0            �R@������������������������       �?���U@Y             a@                            @`�]���@�            0p@������������������������       �v�k		@`             b@������������������������       ���ʳ@D            �\@
                           �?J�l�a@�           �@                           @&21P@           z@������������������������       �_6����@7             X@������������������������       ����rb @�            t@                          �9@��W4B@�             v@������������������������       ���B,3@�            �r@������������������������       �~�a;�@             L@                           �?
�OZ��@�           ޤ@                           @o�q|��	@�            �@                           �?>&���K	@�           `�@������������������������       ����@�            @w@������������������������       �?��Ǣ�	@�           ��@                           �?S+U�=	@[            �b@������������������������       ��^}�A�@!            �N@������������������������       �3��/�@:            �U@                           �?C���@�           ��@                           @�]�7!@�           P�@������������������������       �G.A�P@�            �q@������������������������       �~~d��p@           �x@                           �?��4�p@!           (�@������������������������       ��0�S@'            �Q@������������������������       ����m�@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     r@     �@      2@     �H@     P@      Q@     ��@     @l@     ��@     �t@      A@       @     @U@     �f@      @      @     �`@      "@     @z@      G@     �q@      Q@       @       @     �G@     �U@       @      @     �S@      �?      W@      @@     �V@      A@      �?       @      4@      A@       @      @      <@      �?      I@      5@     �D@      $@                              &@                      *@      �?      ;@       @      .@      @               @      4@      7@       @      @      .@              7@      3@      :@      @                      ;@     �J@              �?     �I@              E@      &@     �H@      8@      �?              5@      ;@                      A@              2@      @      >@      $@      �?              @      :@              �?      1@              8@       @      3@      ,@                      C@      X@      �?      �?      L@       @     �t@      ,@     @h@      A@      �?              7@     �C@              �?      ?@      @     �h@      "@     �U@      6@                      "@      @              �?      ,@       @      =@      @      3@      $@                      ,@      @@                      1@      @     @e@      @      Q@      (@                      .@     �L@      �?              9@       @      `@      @     �Z@      (@      �?              .@     �F@      �?              .@      �?     @_@      @     @U@       @                              (@                      $@      �?      @       @      6@      @      �?      2@     �i@     �x@      .@      F@     �v@     �M@     ��@     �f@     ��@     `p@      @@      2@      \@     `c@      &@      8@     �j@     �B@     �a@     @Y@     �d@     `b@      ;@      &@     �X@     ``@      &@      7@     @g@      ?@      `@     �R@     �c@     ``@      5@      �?      :@      L@      �?      &@      K@      @     �S@      ;@     @P@     �E@      @      $@     @R@     �R@      $@      (@     �`@      9@      I@     �G@     @W@      V@      1@      @      *@      8@              �?      :@      @      *@      ;@      "@      0@      @              $@      "@              �?      @       @      @      ,@      @      "@      �?      @      @      .@                      3@      @      $@      *@      @      @      @              W@     �m@      @      4@     @c@      6@     @z@     �S@     w@     �\@      @              F@     �[@      @      (@     �T@      @      d@      9@      f@      L@      @              5@     �L@              @      F@      @      G@      2@     �M@      8@      @              7@      K@      @       @     �C@             �\@      @     �]@      @@                      H@      `@      �?       @     �Q@      .@     @p@      K@      h@     �M@      �?              $@      @              @      "@       @      @      (@      (@      @                      C@     @^@      �?      @      O@      *@     �o@      E@     �f@     �J@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�q�%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��T��A@�	           ��@       	                    �?��(��@t           �@                          �<@��d�0}@�           �@                          �4@�]�?��@           ��@������������������������       ��t��@�            �s@������������������������       ��ʵ/�5@�             r@                           �?���Ñ>@-            �O@������������������������       ������~@%            �I@������������������������       �Z��h W@             (@
                          �9@���_V	@�           ��@                           @�}l��	@�           P�@������������������������       �&�O�@�           �@������������������������       ��J��@\             b@                            @�(ɓct	@�            �u@������������������������       �dT?>�@�             j@������������������������       �MOCr�@T             a@                            @�%�@K           ��@                           @��U� @�           ��@                           @�7���@�           �@������������������������       ���ICA�@�           ؃@������������������������       �Iؚs @           �x@                           �?	��s�U@           @z@������������������������       �e�A+�@d             c@������������������������       ��2�@@�            �p@                           @\�ޯ[<@�            `q@                           @�%�$�=�?Z            �a@������������������������       ����d'�?,             O@������������������������       ���}��k�?.             T@                           �?����@X             a@������������������������       ��l�,H��?$            �L@������������������������       �D@ӻ�@4            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     @s@     ��@      =@     �M@     �z@     �U@     ��@     �k@     `�@     0w@      4@      .@     �j@     `t@      8@      E@     @s@     �P@     `w@      g@     �w@      n@      1@      �?      R@     @U@      �?      "@     @U@      @     �e@      B@     �b@      I@      @      �?     �P@     @S@      �?      @     �R@      @      e@      =@     �a@     �@@       @              *@     �A@               @     �E@       @     �X@      2@      T@      8@      �?      �?     �J@      E@      �?      @      @@      @     �Q@      &@     �N@      "@      �?              @       @               @      $@              @      @      @      1@       @              @       @               @      @               @      @      @      1@                                                      @               @      @       @               @      ,@     �a@      n@      7@     �@@     �k@     �N@     @i@     �b@     �l@     �g@      *@      $@      Z@     �h@      6@      ;@      g@      <@     `d@     �Z@      f@     �a@      $@       @     @V@     `d@      6@      9@     �c@      3@     �b@     @W@     `d@     @`@      @       @      .@      A@               @      :@      "@      (@      ,@      *@      *@      @      @      B@      F@      �?      @      C@     �@@     �C@     �D@      J@      H@      @              2@      2@              @      =@      9@      4@      >@     �@@      <@       @      @      2@      :@      �?              "@       @      3@      &@      3@      4@      �?      �?      X@      o@      @      1@     �]@      4@     0�@      C@     @y@     @`@      @      �?     @U@     �l@      @      *@     �X@      ,@     ��@     �A@     �t@      \@      �?      �?      N@      d@      �?      @      K@       @     `z@      ,@     �l@     @R@              �?     �F@     �W@      �?      �?      D@       @     `l@      &@     �b@      M@                      .@     �P@              @      ,@             `h@      @     �T@      .@                      9@     @Q@       @       @      F@      @      [@      5@     @X@     �C@      �?              @     �@@       @              "@              J@      @     �@@      &@                      3@      B@               @     �A@      @      L@      ,@      P@      <@      �?              &@      4@       @      @      4@      @      ]@      @      S@      2@       @              @      (@                      ,@      �?     @P@              F@               @              �?      $@                      �?      �?      <@              5@                              @       @                      *@             �B@              7@               @              @       @       @      @      @      @     �I@      @      @@      2@                      �?                       @      @              ?@      @      .@       @                      @       @       @       @      @      @      4@              1@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-�7hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�>fp<@�	           ��@       	                    �?�y��v@}           ܜ@                          �2@E���R�@t           @�@                           �?']T@��@�            t@������������������������       �B�T@]            �a@������������������������       ��4��kL@j            @f@                           @�"+��@�            pp@������������������������       ����i�@�            �m@������������������������       �ϓ(aec@             8@
                           @�[��@	           ��@                           @�J02p~@�           ��@������������������������       ��Bsk[�@�            q@������������������������       �D� ��@7           ،@                            �?�D��L2@+            �P@������������������������       �4`��Z@            �E@������������������������       �Γ(aec@             8@                          �<@��ˊK�@I           $�@                           �?,�m�i>@{           �@                            �?=^sҖ�	@           ��@������������������������       ��)Z�	@           {@������������������������       ������@�             v@                          �7@RU��=@l           ��@������������������������       �;����@V           X�@������������������������       ��mw�@           pz@                           �?�u�x��@�            �t@                           �?*j�bx@8             U@������������������������       ��,�1>@&             K@������������������������       �c�C5@             >@                            �?ֽn���@�             o@������������������������       ��	S��@L            �a@������������������������       ��JQNJ�@J            @[@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     �@      <@      L@     0|@      U@     0�@     �l@     0�@      v@      ?@              Y@     �o@      @      .@      f@      1@     ��@     �V@     Pz@     �`@      $@             �L@     �Q@      @      @     �V@      (@     @\@      M@     �Z@      N@      "@              @@     �H@               @     �L@       @      R@      6@     �I@     �@@      �?              .@      4@                      ;@       @      C@      *@      ,@      ,@                      1@      =@               @      >@              A@      "@     �B@      3@      �?              9@      5@      @      @     �@@      $@     �D@      B@      L@      ;@       @              6@      5@      @      @      9@      $@     �D@     �@@      K@      6@      @              @                               @                      @       @      @      @             �E@     �f@      @      $@     �U@      @      �@     �@@     �s@     @R@      �?              D@     �e@      @      $@     @T@      @     �~@      :@     0s@     �L@      �?              @     �E@      �?      @      C@             �W@      (@      P@      *@                     �A@     @`@      @      @     �E@      @     �x@      ,@     `n@      F@      �?              @      "@                      @      �?      3@      @      @      0@                              @                      �?      �?      *@      @       @      ,@                      @       @                      @              @       @      @       @              ,@      g@     `r@      5@     �D@     0q@     �P@     Pw@     @a@     z@     �k@      5@      &@     �c@     �n@      .@      @@     @m@     �I@     �u@     �Y@     �v@     `c@      4@      $@     �W@     �]@      &@      7@     �^@      =@     �X@     �P@     �^@      S@      ,@      @     �H@     �N@      @      3@      P@      1@     �F@     �I@     �R@      A@      @      @      G@      M@      @      @      M@      (@     �J@      0@     �H@      E@      "@      �?     �O@     �_@      @      "@      \@      6@     @o@      B@     �m@     �S@      @             �A@      U@      @      @     @R@      0@     @c@      "@     �Z@      ?@      @      �?      <@     �E@              @     �C@      @      X@      ;@     ``@      H@              @      :@      H@      @      "@     �D@      0@      9@     �A@     �L@     �P@      �?              @      2@              @      @              (@       @      *@      2@                      @      1@              @      @               @       @      @      0@                              �?                      @              $@      @       @       @              @      7@      >@      @      @     �A@      0@      *@      ;@      F@      H@      �?       @      @      *@               @      3@      (@      @      4@      @@      <@      �?      �?      1@      1@      @      �?      0@      @       @      @      (@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�fvhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?S���mi@�	           ��@       	                    �?3��SX�@"           ܒ@                          �4@����ҷ@B           ~@                          �1@$t��@�            �h@������������������������       �z�ͮ�@0            @R@������������������������       ���͘�l@W            @_@                           �?���a�!@�            �q@������������������������       �yoI�2O@]            �`@������������������������       �:���2�@^            �b@
                            @%�/ƅ@�           ��@                           �?{���@�           ��@������������������������       �|��
��@�            t@������������������������       �*��6��@�            @q@                           @6(��6�?S             `@������������������������       �Pj�K�a @%            �M@������������������������       ��KT^���?.            �Q@                           @��)�E@�           $�@                           �?|�{�~	@�            �@                           @>��fi�	@�           ��@������������������������       ������|	@{           ��@������������������������       ��)�3	@W            �a@                           �?R��D@           �y@������������������������       �\�ڝ�H@[            @b@������������������������       ����,��@�            `p@                            @�t�j�@�           H�@                          �4@���D@]           @�@������������������������       �Y���@.           �}@������������������������       ���䏋@/           �~@                           @v���@z            @i@������������������������       �~4���D@r            �g@������������������������       �lofON@             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      s@      �@      :@      L@     �|@     �U@     (�@     @l@     ��@     0w@     �@@      @     �V@     �c@      @      @     �W@      @     �z@      E@     �r@     @Q@      @      @     �I@     �Q@      @      @      H@       @     @^@      <@     �[@      A@      @              @      >@                      1@       @     @P@      1@      F@      .@      �?              �?      .@                      "@              >@      @      (@      @                      @      .@                       @       @     �A@      ,@      @@      (@      �?      @      F@     �D@      @      @      ?@              L@      &@     �P@      3@       @      @      1@      2@      @      @      .@              <@      @      8@      *@                      ;@      7@                      0@              <@      @      E@      @       @              D@     @U@      �?      �?      G@      @      s@      ,@     �g@     �A@      @              @@      T@      �?             �B@      @     �l@      (@     �d@      ?@      @              1@      G@                      5@      @     �`@      "@     @R@      1@                      .@      A@      �?              0@       @      X@      @     �V@      ,@      @               @      @              �?      "@             @R@       @      ;@      @                      @      @                      @              ;@              0@       @                      @                      �?      @              G@       @      &@       @              1@     �j@     �v@      5@     �H@     �v@      T@     ��@      g@     �@     �r@      :@      1@     �b@      l@      .@      C@     �n@     @P@     @e@      c@     �m@     �h@      6@      1@     �^@     `d@      .@      <@      g@      H@     �Z@     �[@      d@      c@      4@       @     �\@     �a@      .@      9@     �c@      D@      X@     @T@     �c@     `a@      .@      "@      "@      4@              @      <@       @      &@      >@      @      *@      @              <@     �N@              $@      O@      1@     �O@      E@     �S@      F@       @              @      :@               @      =@      @      (@      *@      >@      5@       @              6@     �A@               @     �@@      (@     �I@      =@     �H@      7@                      P@      a@      @      &@     �]@      .@      w@      ?@     @s@     �Z@      @              K@      _@      @      "@     �X@      ,@     `r@      =@      o@     �V@      @              .@     �N@      @      @      <@              f@      0@     �`@      B@                     �C@     �O@       @      @     �Q@      ,@     @]@      *@     @\@      K@      @              $@      (@      �?       @      5@      �?      S@       @      N@      0@      �?              @      "@      �?       @      3@      �?     �R@       @     �M@      0@                      @      @                       @              �?              �?              �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�$�JhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @kw�\@�	           ��@       	                    �?C�����@w           h�@                           �?���@�           �@                            �?���s�@�            �q@������������������������       �����l@l             e@������������������������       �R�L��@M            �[@                            �?�W#�{@�            �v@������������������������       ��J��n�@y            �g@������������������������       ��<��H�@e            `e@
                          �5@K�Ӗf`	@�           ̘@                           �?R!z�#X@�           ��@������������������������       �B����@P           X�@������������������������       ��m�@�            �m@                          �:@�$���	@�           ؉@������������������������       ��\K�r	@J           ��@������������������������       ���Ӧj	@�            �r@                          �4@�H�-�@+           T�@                           @+Ü�@4           0�@                          �1@�Ba�6@�            �m@������������������������       ������?;            @X@������������������������       ��Ц�6�@Y            �a@                          �1@0t��@�           ��@������������������������       �q��á @�            0p@������������������������       �����x@            @y@                           �?��4��@�           x�@                           @�I���@�             y@������������������������       �7P��g@8            �U@������������������������       �/�g��c@�            �s@                          �<@K�؝-@�            �w@������������������������       ��F`��@�            �t@������������������������       �-_دń@'             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     h�@      4@      P@     �}@     @W@     ��@     `j@     �@     0v@      D@      *@     �j@     pt@      ,@     �I@     �t@     �P@     Pw@      e@     0w@     `p@      A@      �?     �L@      X@              &@     @S@       @     �c@      8@     `a@     @Q@      "@      �?      5@      F@              $@      E@       @     �R@      .@     �C@      @@              �?      .@      8@              @      8@              H@       @      3@      8@                      @      4@              @      2@       @      :@      @      4@       @                      B@      J@              �?     �A@             �T@      "@      Y@     �B@      "@              5@      5@              �?       @              E@      @     �O@      6@      "@              .@      ?@                      ;@              D@      @     �B@      .@              (@     �c@     �l@      ,@      D@      p@     @P@      k@      b@      m@      h@      9@      @     �I@      X@      @      0@     �^@      5@     �a@     �P@      b@     �U@      @      @      F@      M@      @      ,@      X@      2@     �S@     �D@     @W@     �P@      @              @      C@      �?       @      ;@      @      O@      9@     �I@      5@              @     @Z@     �`@      "@      8@     �`@      F@     @S@     �S@      V@     �Z@      3@      �?     �Q@     �Z@      @      2@     �S@      9@     �I@     �I@     @P@      G@      .@      @     �A@      =@      @      @     �L@      3@      :@      ;@      7@      N@      @      �?     �R@     �l@      @      *@      b@      :@     P�@     �E@     �z@     @W@      @              :@     @_@       @      @     �J@      @     `y@      0@     `k@      D@      �?              0@     �D@                      (@      @      X@      @     �H@      ,@                      @       @                       @              K@       @      7@      @                      *@     �@@                      $@      @      E@      @      :@      "@                      $@      U@       @      @     �D@      �?     `s@      &@     @e@      :@      �?              @     �@@               @      1@             �a@      @     �G@      &@      �?              @     �I@       @      @      8@      �?      e@       @     �^@      .@              �?      H@     @Z@      @      @     �V@      3@     �j@      ;@     �j@     �J@      @      �?     �@@      P@              @      F@      "@     �[@      "@     �W@      8@      @      �?       @      (@              �?      $@      @      ;@              .@      @       @              9@      J@              @      A@       @      U@      "@      T@      4@      @              .@     �D@      @      �?     �G@      $@     @Y@      2@     @]@      =@                      $@     �A@      @      �?      @@      $@      X@      0@     �Z@      5@                      @      @      �?              .@              @       @      $@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�,]*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�&o��>@�	           ��@       	                   �4@i���@�           Х@                           @R�t�Y@<           ��@                          �0@a$�@G           P�@������������������������       ����@(            �P@������������������������       �����{(@           p|@                           �?]�T=��@�            �@������������������������       ���w8�#�?�            �q@������������������������       ���i�k�@F           H�@
                          �8@Z���n@�           �@                           �?�
��@           ��@������������������������       ��"]�@�            �q@������������������������       �c>�@O           ��@                           �?��w���@�           8�@������������������������       �� �-	@�            �s@������������������������       ��X�-@�            �t@                          �2@R,�}K�@�           ��@                           �?rxV�P@�            �r@                           @.#*̤�@F            �]@������������������������       �� k�ۈ@+            @R@������������������������       ��֤α��?            �F@                           �?�?��Y@k            @f@������������������������       ������@=            �W@������������������������       �,�yl@.            �T@                           �?"<��@           ȉ@                           @5��9�	@�            Pv@������������������������       �9�<d�	@�            `q@������������������������       ��	x���@1            �S@                          �:@1QF�b\@.           @}@������������������������       ��d�!�@�             w@������������������������       �llt�@F             Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     ps@     ��@      7@     �J@     �{@     �R@      �@      k@     h�@     �v@      D@      @      l@     �z@      (@     �A@     @s@     �I@     ؇@     �a@     H�@      n@      =@      �?      Q@     `i@      �?      "@     �^@      *@     �~@     �A@     �q@     �V@      $@      �?     �A@     �S@               @      T@      &@      `@      9@      Y@     �J@       @              @      0@                      @              >@               @      @              �?      @@      O@               @     �R@      &@     �X@      9@      W@     �H@       @             �@@     @_@      �?      @     �E@       @     �v@      $@     �f@      C@       @              "@     �B@                      "@             �d@      @      H@      "@       @              8@      V@      �?      @      A@       @     �h@      @     �`@      =@              @     �c@      l@      &@      :@      g@      C@     �p@     @Z@     q@     �b@      3@       @     @V@     �`@      @      (@      Y@      8@      g@      D@      c@     �N@      &@       @      >@      E@      @      @      =@      @     �U@      @      N@      &@      @             �M@     @W@      @      @     �Q@      2@     �X@     �@@     @W@      I@       @      @      Q@     �V@      @      ,@     @U@      ,@     �U@     @P@      ^@     @V@       @      @     �E@     �G@      @      @     �H@      "@      3@      D@     �C@     �J@      @              9@     �E@      �?      @      B@      @     �P@      9@     @T@      B@       @      "@     �U@     �a@      &@      2@     @a@      7@     Pp@      S@     �l@      ^@      &@              &@      A@      �?      @      =@      @     �Z@      &@      R@      8@                      @      $@                      @       @      M@      @      :@       @                      @      "@                      @       @      ;@      @      ,@       @                              �?                      �?              ?@              (@                              @      8@      �?      @      8@       @     �H@       @      G@      0@                      @      *@      �?      �?      3@       @      *@       @      ;@      ,@                       @      &@               @      @              B@      @      3@       @              "@     �R@     �Z@      $@      .@     @[@      3@     @c@     @P@     �c@      X@      &@      @      @@     �C@      @      (@      I@      &@     �P@      8@     @P@      G@       @      @      @@     �@@      @      $@     �G@      $@     �@@      6@     �G@     �@@       @                      @      �?       @      @      �?     �@@       @      2@      *@              @     �E@     �P@      @      @     �M@       @      V@     �D@     �V@      I@      "@      @      =@     �J@       @      �?     �H@      @     �Q@      6@     �U@     �A@      "@      �?      ,@      ,@       @       @      $@      �?      1@      3@      @      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ0=:+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�y�@M@�	           ��@       	                   �5@�<^��@e           ^�@                           �?��H{r�@�           h�@                           �?��
@�           ��@������������������������       ���;y�e@�            pq@������������������������       ���-��@&           �~@                          �1@5a�ox@�            �u@������������������������       �D	�os @=            @Y@������������������������       �W7���@�            �n@
                           �?!r����	@�           T�@                          �:@���?
@           �@������������������������       ����c	@K           �@������������������������       ��)�U'
@�             t@                            �? FԒ'@�             q@������������������������       �S���@Y            �c@������������������������       �I>���4@H            �]@                          �7@�����@B           h�@                           �?�3)@B           L�@                            �?`����?(           �|@������������������������       ���Ɖ���?B            @Y@������������������������       � �}FN0@�            �v@                           @.�u&B@            �@������������������������       �� ���@           ��@������������������������       ��IOa�@	             4@                            @,R��[�@            px@                          �?@X�eg��@�            @s@������������������������       �iz,U�@�            �r@������������������������       �
4%'V�?             (@                          �9@2���0�@6            �T@������������������������       ��mj � @             C@������������������������       �V�஭@            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     �@      B@      L@      ~@      R@     $�@      m@     ��@     �v@      9@      4@      j@     @s@      ;@     �G@     `s@     @P@     px@     �g@      x@     `o@      3@      "@     @P@     `c@      "@      (@      d@      5@     �n@     �T@     �l@     @^@      @      "@      I@      X@      @       @     �^@      3@     �a@     �J@     �c@     �X@      @      �?      *@     �G@      �?      @      =@      �?     @P@      (@     �S@      =@               @     �B@     �H@      @      @     �W@      2@      S@     �D@      T@     @Q@      @              .@     �M@       @      @     �B@       @     @Z@      =@     �Q@      7@                      �?      1@                      @             �E@      0@      ,@      @                      ,@      E@       @      @      ?@       @      O@      *@     �L@      3@              &@      b@      c@      2@     �A@     �b@      F@      b@      [@     �c@     @`@      ,@      &@      [@     �]@      2@      <@      _@      A@     �W@     �T@     @Z@     �X@      (@             �Q@     �T@      $@      1@     @T@      3@     �P@     �I@     @Q@     �B@      $@      &@      C@     �B@       @      &@     �E@      .@      ;@      @@      B@      O@       @              B@      A@              @      :@      $@     �I@      9@      J@      ?@       @              0@      (@              @      1@       @      =@      3@      @@      ,@       @              4@      6@                      "@       @      6@      @      4@      1@              �?      V@     @i@      "@      "@     @e@      @     �@     �E@      y@     �[@      @              M@      e@       @      @     �Z@      @     �@      6@     �r@     @T@      @              2@     �J@              �?      =@      �?      p@      @     �T@      ,@                              @                       @             @S@              *@       @                      2@      G@              �?      ;@      �?     �f@      @     @Q@      (@                      D@     �\@       @      @     @S@      @     �q@      .@     @k@     �P@      @              D@     @\@      @      @     �Q@      @     �q@      .@     �j@     �P@      @                       @      @              @              @              @                      �?      >@      A@      �?      @      P@             @Y@      5@     �Y@      >@       @      �?      <@     �@@               @     �J@             @Q@      1@     �S@      8@       @      �?      6@     �@@               @     �J@              Q@      1@     �R@      7@       @              @                                              �?              @      �?                       @      �?      �?      @      &@              @@      @      7@      @                       @      �?                       @              3@      �?      @       @                                      �?      @      @              *@      @      2@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJp�.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@��Ҿ6@�	           ��@       	                   �1@lYBo�4@~           ��@                            �?W?�D_@�           ��@                           @jm����@�            �u@������������������������       �� �3`@\             b@������������������������       ���A6j @y            @i@                            @)L���@�            @r@������������������������       ��v6P @U            �`@������������������������       �-Òx�@d             d@
                            @�҅�@�           ��@                           �?C���@           (�@������������������������       ��$���`@�            �j@������������������������       ��(��5�@�           x�@                           @u���@�            �u@������������������������       �ԫ5��!@�             s@������������������������       �)*�@             F@                           �?�#�i@           R�@                           �?��Y�	@t           h�@                            �?�sD�j@�            p@������������������������       �>���7#@`             b@������������������������       ��<3h�@H            @\@                          �:@�?� n�	@�           `�@������������������������       ��F�eZ	@7           0�@������������������������       �N6ɸ�	@�            �l@                           �?��7�'`@�           �@                           �?�/��6@J           ��@������������������������       �m�9\@k            `f@������������������������       ��m5@�             v@                            �?�m� @_           H�@������������������������       �K��7'@U            @_@������������������������       ��U}D!e@
           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     ��@      A@      M@      }@      R@     p�@     �i@     ��@     �u@      ?@       @     @W@      p@      .@      3@     �d@      *@     P�@     @T@     z@     �`@      $@      �?      6@      Z@       @      @     �F@              p@      2@     @a@      G@       @      �?      @     �O@               @      2@             �`@      $@     @S@      B@              �?      @     �C@                       @             �@@      @      ?@      4@                      �?      8@               @      $@              Y@      @      G@      0@                      .@     �D@       @      �?      ;@             @_@       @     �N@      $@       @               @      .@                      0@              O@       @     �@@               @              *@      :@       @      �?      &@             �O@      @      <@      $@              �?     �Q@     @c@      *@      0@      ^@      *@     �v@     �O@     pq@     �U@       @              F@     �]@      $@       @      T@      @     0q@     �E@     �f@     �P@      @              1@      <@      @      �?     �@@       @      >@      <@      B@      =@      @              ;@     �V@      @      @     �G@      @     �n@      .@     @b@     �B@              �?      ;@     �A@      @       @      D@       @     @U@      4@     @X@      5@      @      �?      ;@      ?@      @      @      A@      @     �S@      &@      V@      2@      �?                      @               @      @      @      @      "@      "@      @       @      .@      h@     �s@      3@     �C@     �r@     �M@     @x@      _@      y@     @k@      5@      .@     @^@     �d@      0@      ;@     �d@     �@@     @Z@     �S@     �a@     �^@      ,@             �E@      K@       @      &@      9@              <@      .@     �H@      <@       @              ;@      =@      �?      @      ,@              &@      @      :@      7@       @              0@      9@      �?      @      &@              1@      "@      7@      @              .@     �S@     @\@      ,@      0@     �a@     �@@     @S@     �O@     @W@     �W@      (@      @      M@      U@      "@      $@     �Y@      *@      K@     �H@     �Q@     �I@      &@       @      4@      =@      @      @      C@      4@      7@      ,@      7@     �E@      �?              R@     `b@      @      (@     �`@      :@     �q@      G@      p@      X@      @              ?@     �S@      �?      (@     �N@      &@     @c@      *@     �\@      H@      @               @      ?@                      .@      @     @T@      @      >@      @                      7@      H@      �?      (@      G@      @     @R@      $@     @U@      E@      @             �D@      Q@       @             @R@      .@      `@     �@@     �a@      H@      �?              0@      &@      �?              2@      "@     �A@      @      2@      $@      �?              9@     �L@      �?             �K@      @     �W@      ;@     @_@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�*�/��@�	           ��@       	                    �?�5� ��@�           ��@                            �?�DΕ@�           Ȅ@                           �?��H*�@�             j@������������������������       �0�1+G2@^            �b@������������������������       �ɇ��b@$            �M@                           �?u� Ѷ@"           �|@������������������������       ��؞m.@�            �m@������������������������       ��iA�E�@�            �k@
                           �?>��#��	@�           ̘@                           �?MWyXi�	@�           ԑ@������������������������       ��s7=.i@�            �y@������������������������       ���s��p
@�           �@                            �?�O�:�@           �{@������������������������       �xe��|o@T            �`@������������������������       �h�D�,@�            �s@                           �?C�A"N@8           ��@                          �4@�Wro� @m           ��@                           @�WD-*�?�            �u@������������������������       �V���k��?�             m@������������������������       �v��6�@A            �\@                          �5@�+�dc@�            �k@������������������������       ����'Ο @"            �H@������������������������       ��|F�Ia@k            �e@                          �7@d�H [�@�           �@                           @ �� �w@
           ��@������������������������       �ӭ�S1�@�           ��@������������������������       �����
Y@|             h@                            @���3�@�            �r@������������������������       ������@�            �n@������������������������       ��Y]g@&            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        =@     �q@     ��@     �E@     �O@     |@     @R@     ��@     �k@     �@     �x@      8@      ;@     `g@      u@     �@@      G@     �s@     �N@     @z@     @g@     �u@      q@      5@       @      M@      W@      @       @      V@      @     �f@      @@     ``@      O@      @       @      *@      A@               @      6@      @     �M@      @     �F@      6@               @      &@      ?@              �?      1@      �?     �A@      @      <@      1@                       @      @              �?      @       @      8@              1@      @                     �F@      M@      @      @     �P@      @     @^@      :@     �U@      D@      @              7@      7@      @      @      @@       @     �Q@      .@     �@@      >@      �?              6@     �A@              �?      A@      �?     �I@      &@     �J@      $@       @      9@      `@     �n@      >@      C@     `l@     �K@      n@     @c@     �j@     �j@      2@      9@     �Y@     @e@      :@      :@      e@     �D@      a@     @Z@     �c@     �d@      1@      @      5@     @S@      @      @     �O@       @     @Q@     �A@      M@      L@      @      6@     @T@     @W@      3@      3@     �Z@     �@@      Q@     �Q@     @Y@      [@      *@              ;@      S@      @      (@      M@      ,@     �Y@     �H@      K@      H@      �?              @      7@              �?      8@      @      C@      *@      "@      *@      �?              6@     �J@      @      &@      A@       @     @P@      B@     �F@     �A@               @     @W@     @m@      $@      1@     �`@      (@     Ђ@     �B@     �x@     �^@      @              (@     @Q@      �?      �?      A@             Pq@      @     �`@      A@      �?              @     �@@              �?      .@              h@       @     �S@      0@      �?              @      3@                      @             �a@      �?     �J@      @                      �?      ,@              �?      "@             �I@      �?      :@      $@      �?              @      B@      �?              3@              U@      @     �K@      2@                      �?      "@                       @              5@      �?      "@                              @      ;@      �?              &@             �O@       @      G@      2@               @     @T@     �d@      "@      0@      Y@      (@     Pt@      @@     Pp@      V@       @             �H@     �_@      @       @     �J@      "@     �p@      ,@     `h@     �N@       @             �B@     �X@       @       @     �B@      @      k@      (@     `b@      C@      �?              (@      <@      @      @      0@      @      I@       @      H@      7@      �?       @      @@      C@      @       @     �G@      @      M@      2@     �P@      ;@               @      >@      B@       @      @      F@      @     �B@      0@     �I@      5@                       @       @       @      @      @              5@       @      .@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�I�
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��b��=@�	           ��@       	                   �<@30��@:           ��@                           �?fj6��@�           ��@                           �?|)RcH�@w           �@������������������������       �mN�Ė�@            |@������������������������       ��a�VD@j             d@                           @��6�~	@(            �@������������������������       ��"�A]	@           $�@������������������������       ���@��A@            �K@
                            �?�%@�             n@                           �?[W�
�4@I            @\@������������������������       ���r�@>            �W@������������������������       ��J�r�@             2@                           @�> �@R             `@������������������������       ��w�A��@.            �R@������������������������       ��x�k�R@$             K@                            @yFxk�@h           ؛@                          �7@9WH��@�           �@                           @p#,C`@�           ��@������������������������       ���<�@�             p@������������������������       ��b0WO@,           `�@                            �?t,�c�@�            �t@������������������������       ���tN�e@�            �i@������������������������       �P����?@R             `@                           �?+�mE�@�            �s@                           @��%�k{�?M            ``@������������������������       �g�2dj]�?!             K@������������������������       ����=S�?,            @S@                           @O�@�f�@|            @g@������������������������       ���ƄW?@L             \@������������������������       �W��6�V@0            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      s@      @      9@     �L@     �{@     �U@     \�@     �m@     ��@     u@      B@      0@      j@     �r@      1@      E@     �r@     �Q@     0w@     �h@     0w@     �j@      >@      .@     @f@     �p@      0@      B@     �p@      L@     �v@      d@     �u@     �b@      <@      �?      P@     �S@      @      @     �Q@      @     �d@      ;@     `c@      A@      @      �?      G@      Q@      @      @     �L@      @     �[@      :@     �Y@      8@      @              2@      $@                      ,@              K@      �?     �J@      $@              ,@     �\@     �g@      *@      @@     �h@     �I@     �h@     �`@     �h@     @]@      8@      (@      \@     �g@      *@      @@     �g@      H@     �g@     @]@     �g@     �\@      2@       @       @       @                      $@      @      @      1@      @       @      @      �?      ?@      <@      �?      @      =@      ,@      &@      B@      4@      O@       @      �?      @       @              �?      $@      $@      @      2@      "@     �E@       @      �?      @       @                      @      $@      @      .@      @      D@                      @                      �?      @                      @      @      @       @              8@      4@      �?      @      3@      @      @      2@      &@      3@                      &@      (@      �?      �?       @       @      �?      2@       @      (@                      *@       @              @      &@       @      @              @      @                     @X@     @i@       @      .@     @b@      0@      �@     �C@     P|@      _@      @             �U@     �f@      @      *@     �\@      *@     ��@     �@@      w@     �Z@      @             �M@     �b@      @      $@     �Q@      "@     �}@      7@     0p@     @Q@      @              4@      B@       @              0@       @      X@      $@      H@      3@      �?             �C@      \@      �?      $@     �K@      �?     �w@      *@     `j@      I@       @              <@     �@@      �?      @      F@      @      O@      $@     @[@     �B@       @              3@      6@               @      3@      @     �B@      @     �P@      =@                      "@      &@      �?      �?      9@      �?      9@      @      E@       @       @              $@      5@      @       @      ?@      @      a@      @     @U@      2@      �?              @      @                      @       @     @R@      @     �@@      @                       @      @                               @      A@       @      &@                              @                              @             �C@      @      6@      @                      @      2@      @       @      ;@      �?     �O@              J@      *@      �?              �?      ,@              �?      3@              C@             �A@      @                      @      @      @      �?       @      �?      9@              1@      "@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��'6pF@�	           ��@       	                   �5@!��f�@|           P�@                           �?�����`@�           ��@                          �2@Na\�@�             v@������������������������       �yq�5h@l            @e@������������������������       ����4�@x             g@                           @�I���-@�           �@������������������������       �u�vB��@K           H�@������������������������       �����U@�             o@
                          �<@b�����	@�           �@                           �?��Ay�	@%           �@������������������������       ��u �d�	@�           P�@������������������������       �ޫ�Τ�@�             k@                           @ے�� 		@�             l@������������������������       �������@�            @i@������������������������       ��w�Z@             7@                            �?z (�/?@8           ��@                           @4`&I<@           �z@                           @���y��@K            �_@������������������������       �`��� @;             X@������������������������       �C{T5�j@             ?@                           �?�<�C]@�            �r@������������������������       �܉W�h@_             d@������������������������       ��x�#� @X            �a@                          �<@�'�d�@6           Г@                           @�=��j@           �@������������������������       ��I�>@           8�@������������������������       �)#v���@�            0w@                          �=@]�E�M@'             M@������������������������       ��}W�J�?             .@������������������������       �~<R*�@            �E@�t�b��
     h�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     `�@      :@      O@     {@     �T@     0�@     `j@     P�@      w@      >@      0@     �j@     �t@      3@     �F@     �r@     @P@     �x@     �d@     �w@     0p@      6@      @     �S@     �e@      @      ,@     `b@      7@      p@     �Q@     `k@     �_@      @              7@     �F@               @      @@             @\@      *@     @V@     �A@       @              @      <@                      5@              K@      @      D@      3@                      3@      1@               @      &@             �M@      "@     �H@      0@       @      @      L@      `@      @      (@     �\@      7@     �a@     �L@     @`@      W@      @      @      A@      T@       @      @     @V@      .@      V@      @@     @X@      R@                      6@      H@       @      @      :@       @     �K@      9@     �@@      4@      @      &@     �`@     �c@      .@      ?@     �c@      E@     �a@      X@      d@     �`@      .@      &@     �Z@     �^@      *@      2@      `@      ?@      `@     �R@     @`@     �V@      *@      &@      T@     @Z@      *@      .@     �W@      ;@     �S@     �L@     �V@     �P@      *@              ;@      1@              @      A@      @     �H@      2@      D@      9@                      <@      B@       @      *@      <@      &@      (@      5@      ?@     �D@       @              8@     �@@       @      *@      :@       @      (@      .@      <@      D@      �?              @      @                       @      @              @      @      �?      �?              Y@      l@      @      1@     @`@      2@      �@     �F@     �x@     @[@       @              8@      H@      �?      �?     �@@      @     �h@      @     @W@      7@                      &@      5@      �?              @             �K@      @      2@      (@                      �?      0@                      @             �G@      �?      .@      &@                      $@      @      �?                               @      @      @      �?                      *@      ;@              �?      <@      @     �a@      @     �R@      &@                      @      .@              �?      5@       @     �P@             �F@      @                      "@      (@                      @      �?     �R@      @      >@      @                      S@      f@      @      0@     @X@      .@     �{@      C@     s@     �U@       @             @Q@     �e@       @      ,@      U@      .@     @{@      C@     �r@     �R@       @             �H@     �]@               @     �H@      (@     0u@      2@      j@      C@      @              4@      L@       @      (@     �A@      @     @X@      4@     �U@      B@      @              @      @      @       @      *@               @              "@      (@                       @                              @              @                      �?                      @      @      @       @      @               @              "@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @1�n,�1@�	           ��@       	                   �<@$�.�U�@k           t�@                           �?�WHh@�           �@                           �?`Y��J@�           Ȉ@������������������������       ���-�@�            �q@������������������������       ��{����@;           �@                           �?���I@�           ��@������������������������       �ɢ���@           ؊@������������������������       �׹+���@�            u@
                           �?�N���	@�            �n@                           �?U�5-�@%             M@������������������������       �b �K:�@
             3@������������������������       ����%ԭ@            �C@                            �?�:8	@~            `g@������������������������       �O_ ���@B            �Y@������������������������       �n��D�^	@<            @U@                            �?�e7��@           <�@                           @�b�Aa?@�            �w@                          �5@��.+ϟ@�            pu@������������������������       �J�
>�W�?�            �m@������������������������       ���h7@I            �Z@                          �4@+&#���@            �@@������������������������       �8�&2 @	             1@������������������������       ���b}@
             0@                           @Y�����@)           \�@                           @����K@�           h�@������������������������       ���
��@�           ��@������������������������       ���˅E�?             .@                           �?~c��b@{           P�@������������������������       ��-���(@�            �s@������������������������       ����Z@�            �r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@      p@     ��@      ?@      L@      z@      Q@     �@      l@     0�@      x@      D@      ,@     �g@     �v@      4@     �E@      r@      K@     �x@      g@     �w@     `p@     �A@      &@     �d@      u@      0@      C@     Pp@      C@     �w@     �b@     Pv@     �i@      A@              M@     �a@      "@      (@     �X@      2@     �d@     �P@     @[@     �X@      0@              3@      C@      @       @      B@      @     �X@      &@      E@      9@                     �C@     @Z@      @      @     �O@      .@     @P@      L@     �P@     @R@      0@      &@     �Z@      h@      @      :@     @d@      4@     �j@     �T@      o@     �Z@      2@      &@     @U@     �_@      @      9@     �^@      *@     �`@     �N@     �e@     �T@      2@              6@     �P@      �?      �?      D@      @      T@      6@     �R@      8@              @      8@      =@      @      @      ;@      0@      5@      A@      8@     �L@      �?              @       @              �?      &@              "@       @      @      (@      �?              @       @                      @              @                      @                              @              �?      @              @       @      @      "@      �?      @      4@      5@      @      @      0@      0@      (@      :@      4@     �F@              �?      @      "@               @      @      $@      @      6@      ,@      <@               @      *@      (@      @       @      *@      @      @      @      @      1@                     @Q@     �l@      &@      *@      `@      ,@     p�@      D@     �|@     �^@      @              9@     �A@      @              ;@      @      e@      *@      R@      =@                      6@     �@@       @              ;@      @     �c@       @     �Q@      5@                      @      7@                      0@             �^@      @      L@      &@                      2@      $@       @              &@      @      A@      @      ,@      $@                      @       @       @                              &@      @       @       @                               @                                      @       @      �?      @                      @               @                              @      @      �?      �?                      F@     `h@      @      *@     @Y@      &@     `z@      ;@     x@     @W@      @              <@     �Q@       @      �?      K@      "@     @p@      ,@     @i@     �D@      @              <@     �Q@       @      �?     �G@      @     @p@      &@     @i@     �C@      @                                              @      @              @               @                      0@      _@      @      (@     �G@       @     @d@      *@     �f@      J@       @              "@     �P@      @       @      :@      �?     @V@      �?     �T@      :@                      @     �L@              @      5@      �?     @R@      (@      Y@      :@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ]��%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Vl<�6@�	           ��@       	                    �?��[n�@           �@                          �5@��LX�@/           �~@                           �?4�5�@�            �p@������������������������       ��W��6�@E            @\@������������������������       �V�~��@X            �b@                           �?h�+�l@�            @l@������������������������       ��5���@/             R@������������������������       �]1/fpl@c            @c@
                            �?�c���@�           ��@                          �8@��x�@s            `g@������������������������       �Ë�����?g            �d@������������������������       ��7�g�@             6@                           @���1��@_           �@������������������������       ��%@Sz@�            Pu@������������������������       ���U��@�            �i@                            @$��@�           �@                          �1@��X�=�@�           d�@                           @c�PW@�            �q@������������������������       ��gɓ�@F            @[@������������������������       ���Bn�: @t            @f@                           �?[ե.n@�           �@������������������������       ���w�<�@E            @[@������������������������       �-c�9�@�           4�@                          �1@y�ߊ�@�           P�@                           �?���:�@7            �S@������������������������       ����� @             1@������������������������       ���Z^�l@+             O@                           @�L3�z	@�           ؆@������������������������       ���~� �	@V           ��@������������������������       �����@^            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     Pq@     0�@      @@     �G@     �~@     �Q@     ��@      j@     ��@     0v@     �C@      �?     @S@      e@      �?      $@     �Z@      @     `{@      I@     �q@      S@      @      �?      J@     @S@              "@      L@      �?     �Z@      ?@     @Z@     �G@      @              :@      B@              @      3@      �?     �S@      .@     �O@      3@      @              "@      "@               @      "@      �?      E@      @      6@      $@      @              1@      ;@              �?      $@             �B@      "@     �D@      "@              �?      :@     �D@              @     �B@              ;@      0@      E@      <@       @      �?      @      (@                      .@              (@              *@      &@      �?              3@      =@              @      6@              .@      0@      =@      1@      �?              9@      W@      �?      �?     �I@      @     �t@      3@     �e@      =@      �?              �?      3@      �?              5@      @     @V@      �?     �E@       @      �?              �?      2@      �?              0@             �U@              D@      @                              �?                      @      @      @      �?      @      @      �?              8@     @R@              �?      >@      @     `n@      2@     �`@      5@                      6@      C@                      1@      @      e@      $@     �Q@      *@                       @     �A@              �?      *@             �R@       @      O@       @              3@      i@     �w@      ?@     �B@     �w@     �O@     Ё@     �c@     Ȁ@     pq@     �@@      *@     ``@     �o@      *@      7@     pp@      F@     �{@      \@     �w@      h@      0@      @      "@     �G@              �?      ,@      �?     �\@      "@      O@      8@              @      @      :@                      @      �?      =@      @      0@      *@                       @      5@              �?      "@             �U@       @      G@      &@               @     �^@      j@      *@      6@      o@     �E@     `t@     �Y@     �s@      e@      0@      @      "@      "@              @      ;@      @      @      $@      <@      @       @      @     @\@     �h@      *@      3@     �k@     �B@      t@     @W@     �q@     `d@      ,@      @     @Q@     �_@      2@      ,@     �]@      3@      `@     �G@      d@     �U@      1@              @      2@      �?      �?       @              ?@       @      ,@      @                      @                                              @       @       @       @                       @      2@      �?      �?       @              8@              (@       @              @     �O@      [@      1@      *@     @]@      3@     �X@     �F@     @b@     �T@      1@      @      N@     @X@      *@      &@     �W@      2@     �N@     �D@     @W@      O@      .@              @      &@      @       @      6@      �?     �B@      @     �J@      4@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJr��2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���q@�	           ��@       	                    �?>���m�@g           R�@                          �<@��ɽم@�           Ȅ@                           �?��k��@s           H�@������������������������       ��	�a�@�            q@������������������������       ��y�>L@�            �s@                          �=@���0��@+             T@������������������������       ��y+� @             A@������������������������       ���T�@             G@
                           @�$��m	@�           @�@                           �?c�+z�<	@J           �@������������������������       ������v	@n           P�@������������������������       �:
���@�            �u@                           �?S�GCL	@            �i@������������������������       ��w���@T             a@������������������������       ��Ċ>��@+             Q@                           �?.�鵹@/           ��@                           @a��SI)@n           �@                            �?���9���?�            �x@������������������������       � Dg�ֳ @�            `i@������������������������       �c�����?x            �g@                           �?��l�H@v             g@������������������������       ��mw�U� @=             Y@������������������������       �}RX�@9            @U@                          �3@,���+@�           t�@                            �?�P��9b@           {@������������������������       ��/���?>            �Y@������������������������       ��>�9Q�@�            �t@                          �<@�1��|_@�           `�@������������������������       ��|�Z@�           `�@������������������������       �x]
�@,             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     `s@     ��@      @@      K@     @      T@     ��@      l@      �@     pw@      @@      *@      k@     @r@      8@     �F@     Pv@     �M@     �u@     @h@     �w@     �p@      ;@             �Q@     �X@      �?      @     �S@      @     �b@     �A@      c@     �O@      @              L@     @U@      �?      @     �Q@      @     �a@      ;@     �b@      F@      @              1@     �F@      �?      @      D@      @     @R@      1@     �M@      *@                     �C@      D@                      ?@      �?      Q@      $@     @V@      ?@      @              .@      ,@               @       @               @       @      @      3@       @              @       @                                              @       @      ,@                      "@      @               @       @               @      @       @      @       @      *@     @b@      h@      7@      C@     `q@     �K@     �h@     �c@      l@     `i@      6@      $@     �`@     �c@      6@     �A@      o@      F@     @f@      ^@      j@     `f@      ,@      $@     �X@     @^@      4@      ;@     �h@     �A@     @Z@      W@     `b@     �`@      *@             �@@     �A@       @       @     �H@      "@     @R@      <@      O@     �F@      �?      @      ,@     �B@      �?      @      >@      &@      4@     �C@      .@      8@       @      @      "@      9@      �?              :@      @      $@      7@      @      3@       @              @      (@              @      @      @      $@      0@       @      @               @     @W@     @n@       @      "@     �a@      5@     �@      >@     �z@     @[@      @              3@     @S@      �?              ?@      @     @q@      @     @a@      7@      @              *@      I@                      1@      @     �i@       @     @V@      *@                      @      B@                      $@       @      X@       @      F@      "@                      "@      ,@                      @       @     �[@             �F@      @                      @      ;@      �?              ,@      �?     �Q@      @     �H@      $@      @               @      *@                      $@      �?     �F@              9@      @                      @      ,@      �?              @              9@      @      8@      @      @       @     �R@     �d@      @      "@     @[@      0@     �t@      8@      r@     �U@       @              .@     �Q@      @      �?      9@              c@      @     �`@      :@                       @      .@                      @             �J@      @      7@      @                      *@      L@      @      �?      6@              Y@      @     @[@      7@               @     �M@     �W@      @       @      U@      0@     �f@      2@     �c@      N@       @       @     �G@     �U@       @      @     �P@      0@      f@      2@     @b@     �I@       @              (@      @      �?      �?      2@              @              (@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJp)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@g���H@�	           ��@       	                    �?����@�           x�@                           @�*���@�            �s@                           �?����@�            �o@������������������������       �Q'���f@@            �Z@������������������������       ���X2~@e            @b@                           �?�.�$@*            �P@������������������������       �Q�V#k@             2@������������������������       �U��$@             H@
                           @7H�n�@�           ��@                          �1@{)l�8@h            �e@������������������������       �9.�.��@9             V@������������������������       ��m�@/            @U@                            �?���!@� @_           ��@������������������������       ���W�(@�            u@������������������������       �][�Z��?�             l@                          �<@�uD��@�           V�@                           �?�Lc��@+           ��@                          �9@௭�Ԥ@�           �@������������������������       �j1��^@           8�@������������������������       ���>�}@G            �^@                            @+ͼ�p@e           �@������������������������       �HK�4�@           ��@������������������������       �hϦ�u�@Q           ��@                          �=@8�-�5|	@�             u@                            �?��lׂ�@=             W@������������������������       ���w�U�@#             I@������������������������       �������@             E@                           @��6֍	@�            �n@������������������������       �g�W�*[	@w             h@������������������������       ��
և&*@             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     Pr@     �@      ?@      K@      }@     �T@     ��@      l@     P�@     `v@      7@       @     �F@     `b@      @      "@      T@      @      {@     �D@      i@     @V@               @      6@     �I@      @      �?     �F@      �?      S@      6@     �I@     �F@               @      *@      >@      @             �B@             �P@      2@     �F@      C@               @      @      0@      @              ,@              C@      @      &@      ,@                      $@      ,@                      7@              =@      (@      A@      8@                      "@      5@              �?       @      �?      "@      @      @      @                      �?      @                      @              @                      @                       @      .@              �?      @      �?      @      @      @       @                      7@      X@      �?       @     �A@       @     `v@      3@     �b@      F@                       @      7@              �?      "@      �?     @R@      ,@      @@      2@                       @      (@                       @              A@      "@      4@      "@                              &@              �?      @      �?     �C@      @      (@      "@                      5@     @R@      �?      @      :@      �?     �q@      @     @]@      :@                      @     �E@      �?      @      .@      �?      e@       @     �Q@      6@                      ,@      >@                      &@             @]@      @      G@      @              2@      o@     �z@      ;@     �F@      x@     �S@     �@     �f@     �@     �p@      7@      .@     �j@     �w@      8@     �A@     u@      L@     (�@     `b@     �@      i@      3@      @      O@     �[@      @      @      R@      @     �m@      1@     `g@      @@      �?              K@     @V@      @      @     �I@      @     �i@      ,@     `c@      ?@      �?      @       @      6@                      5@       @      >@      @      @@      �?              (@     �b@     �p@      5@      =@     �p@      I@     �s@     @`@     pv@      e@      2@      "@      W@     �i@       @      ;@      e@      A@      m@     �V@     �p@     �[@      "@      @      M@     �P@      *@       @      X@      0@     �S@      D@     �V@      M@      "@      @      B@      F@      @      $@     �G@      7@      >@      B@      @@      Q@      @      �?      (@      $@      �?      @       @      @      @      @      ,@      ;@              �?      @      @               @       @      @       @      �?      @      7@                       @      @      �?       @      @              @      @      @      @               @      8@      A@       @      @     �C@      3@      8@      ?@      2@     �D@      @       @      4@      <@              @      ;@      0@      .@      >@      (@      @@      @              @      @       @              (@      @      "@      �?      @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�k!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��7Fd@�	           ��@       	                    �?8�x=@           �@                           �?y��ĳ*@�           H�@                            @Ҷ`��@�            �l@������������������������       �x��M�@O            �_@������������������������       ���3o�K@@             Z@                            �?Ļ�Z��@           0z@������������������������       �M��W,3@�            �l@������������������������       ��Z/��� @x            �g@
                           �?��F��@t           �@                            �? <�qL�@�            �m@������������������������       ����L�@O            �^@������������������������       ��<�u4�@G            �\@                          �7@?vP4��@�             u@������������������������       �i��J! @�            0p@������������������������       �ɯ��R@0            @S@                           @�D��^X@�           �@                           �?ᬵ1-w	@�           ؗ@                           @��� Q	@\           ؀@������������������������       �����j�@�            @n@������������������������       ��<>4&�@�            �r@                           @����oe	@o           ؎@������������������������       ��2�X;	@           ؊@������������������������       �TG�>�@P             `@                           @��Q�@�           4�@                           @�G��Ԙ@�           @�@������������������������       ��
Pr�@            �i@������������������������       ����i�@           �@                          �;@A*JS�@V            @_@������������������������       �F1_ @L            �[@������������������������       ��"�@}��?
             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@      t@     �@     �C@     �M@     `}@      R@     X�@     �j@     `�@     @t@      :@              S@      d@      @      *@     �W@      @     �|@     �F@     �q@     �Q@      @             �A@      T@       @      &@      N@      @      q@      =@      ]@      C@      �?              *@      @@       @       @      @@      �?     �P@      5@     �B@      1@      �?              @      3@               @      7@      �?      @@      *@      2@      $@      �?              @      *@       @      @      "@              A@       @      3@      @                      6@      H@              @      <@      @     �i@       @     �S@      5@                      ,@      7@              @      3@      @     �]@      @      ?@      .@                       @      9@                      "@             �U@      @      H@      @                     �D@      T@       @       @     �A@       @     �g@      0@     �d@     �@@      @              >@      G@               @      4@              J@      "@      M@      2@       @              @      9@              �?       @              8@              E@      *@       @              7@      5@              �?      (@              <@      "@      0@      @                      &@      A@       @              .@       @     @a@      @     @[@      .@      @              "@      9@       @              @              _@      @     �S@      "@       @               @      "@                       @       @      ,@      @      ?@      @      �?      9@     �n@     0z@     �A@      G@     pw@     @P@     �@      e@     @     �o@      4@      7@      f@     �o@      <@     �A@     �o@     �F@      f@     �b@     @i@      e@      .@      @     @Q@     �Y@      3@      @     �U@      0@      O@     �G@      N@      N@      @      @      @@     �B@      *@      �?      E@      (@      B@       @      >@      <@              @     �B@     @P@      @      @      F@      @      :@     �C@      >@      @@      @      0@      [@      c@      "@      =@     �d@      =@     �\@     �Y@     �a@     @[@      $@      "@     @V@     @`@      "@      =@     �b@      7@     @Y@      S@      a@      Y@      @      @      3@      6@                      1@      @      *@      :@      @      "@      @       @     @Q@     �d@      @      &@     �^@      4@     �v@      4@     pr@      U@      @       @     �H@      c@      @      $@      [@      1@     �t@      .@      q@     @R@      �?       @      &@      >@      �?      @      ;@      $@     �L@      $@     �D@      *@                      C@     �^@      @      @     @T@      @     Pq@      @     �l@      N@      �?              4@      (@      �?      �?      ,@      @      ?@      @      7@      &@      @              3@      &@      �?      �?      @      @      ?@      @      5@       @      @              �?      �?                       @                               @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��QmhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?`$���k@�	           ��@       	                    �?�>@M	@           H�@                            �?�"*>�@�           ��@                          �4@�6<6��@x            `e@������������������������       �ՄǄ�@0            �O@������������������������       �>��x#2@H             [@                          �=@"�*�%�@           �z@������������������������       �QJw�K@           `x@������������������������       �BR��@            �A@
                           �?�UF���	@�           ��@                           �?M{#���@�            �r@������������������������       ����$�@V            @`@������������������������       �&�I ��@l            �d@                           �?�+h��
@�           ��@������������������������       ��.BV7	@�            �l@������������������������       �1����	@@           �~@                           �?V��&$@�           �@                           �?T��K�K@�           ��@                            �?/2�1�@           �|@������������������������       ����l���??            �X@������������������������       �����Q@�            pv@                          �=@�;�|�#@�            �r@������������������������       �Z�t^7@�            �q@������������������������       �+�%W�@	             0@                           @�n�)@�           �@                           �?	��	!�@�           (�@������������������������       ���m�@�            �o@������������������������       �����@            �z@                          �7@�)4]j2@-            �@������������������������       �~헮}�@�           P�@������������������������       ���4�{@�            �n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     @s@     �@      ?@      L@     �{@     �W@     x�@     �m@     ��@     �u@      ?@      ,@     �e@     �m@      5@      <@     �n@     �N@     �k@     �b@     `p@      f@      8@      @     �C@     �V@      @      "@     �V@      &@     @\@     �D@     �_@     �O@      @      �?      @      *@              @      8@       @      H@      2@      C@      ,@      �?                      @                      @       @      4@      @      6@      @              �?      @      "@              @      4@              <@      (@      0@      "@      �?       @      @@     @S@      @      @     �P@      "@     @P@      7@      V@     �H@      @       @      =@     @S@      �?      @     �O@       @     �O@      3@     �T@     �B@      @              @              @              @      �?       @      @      @      (@              &@     �`@     �b@      0@      3@     �c@      I@     @[@     �[@      a@     �\@      3@              B@     �F@      @      @     �D@      @     �L@      9@      I@      <@       @              *@      .@      @      @      6@      @      9@      &@      5@      &@                      7@      >@              �?      3@              @@      ,@      =@      1@       @      &@     @X@      Z@      *@      (@     �\@     �G@      J@     @U@     �U@     �U@      1@       @      @@     �A@      @              8@      ,@      0@      <@      7@     �F@      @      "@     @P@     @Q@      @      (@     �V@     �@@      B@     �L@     �O@     �D@      &@      �?      a@     @s@      $@      <@     �h@     �@@     ��@      V@     ��@     @e@      @             �A@      W@              @     �G@      $@     �u@      0@     �e@      ;@       @              2@      N@              @     �A@      @     `k@      @     �V@      0@                              "@              �?      @      @      I@              9@      @                      2@     �I@              @      <@      @      e@      @     @P@      *@                      1@      @@                      (@      @     �_@      $@     �T@      &@       @              1@      @@                       @      @     �^@      @     �T@      "@      �?                                              @              @      @      �?       @      �?      �?     @Y@      k@      $@      5@      c@      7@     �{@      R@     Pv@     �a@      @      �?      N@     �Y@      �?      @      P@      0@     `f@     �I@     @_@     �Q@      �?      �?      7@     �@@              @      ;@      @      J@      1@      O@      >@      �?             �B@     @Q@      �?      @     �B@      (@     �_@      A@     �O@      D@                     �D@     �\@      "@      ,@      V@      @     Pp@      5@      m@     @R@      @              >@     �T@      @       @     �J@      @     �j@      @     `e@      F@       @              &@      @@      @      @     �A@      @      G@      0@     �N@      =@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJhw1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @��<�Q@�	           ��@       	                    �?g���@y           ��@                          �;@���J��@�           p�@                           �?C�D��@i           X�@������������������������       ���ضc@           �x@������������������������       �x���@a            �c@                            �?�C�
�@8            �X@������������������������       �E���@            �G@������������������������       �x�	bi�@             J@
                           �?lgW>	@�           ̘@                          �;@��uo&�	@�           D�@������������������������       ����W�	@>           �@������������������������       ���T\-&
@�            �n@                          �3@���١@            z@������������������������       �[���@b             c@������������������������       �m��Z9J@�            �p@                           @�xK9�@$            �@                           �?Q4��@�           $�@                           @��~.��?�            �u@������������������������       ��X�ka @�            `n@������������������������       ����t��?D            �Z@                            @Â����@
           `�@������������������������       ������@�           `�@������������������������       �3a��]��?@             X@                           @,����@<           �@                           @�y,�*Z@5           �~@������������������������       �G�+���@�            �w@������������������������       �	�
to�@F            @]@������������������������       �i	\��p @             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        9@     pq@     ��@      8@      L@      ~@     �R@     Ȏ@     �l@     P�@     @v@      ?@      8@     �g@     �v@      .@     �F@     �u@      K@     @v@      i@      x@     @m@      ;@      �?     �K@     �X@       @      $@     �S@       @     `b@     �B@      d@      M@      @              E@     �U@       @       @     �N@       @     �a@      :@     �a@     �D@      @              @@     @Q@       @       @      H@             �W@      6@     �V@      =@      @              $@      1@                      *@       @     �H@      @     �H@      (@              �?      *@      (@               @      1@              @      &@      5@      1@      �?      �?      @      @                      @                      @       @      .@      �?              @      "@               @      (@              @      @      *@       @              7@     �`@     �p@      *@     �A@     �p@      J@      j@     �d@     �k@      f@      6@      7@     �[@     �h@      *@      ;@     �j@     �D@      _@     �\@     @c@     �`@      3@       @      U@      c@      &@      1@     `g@      ;@     �Z@     �W@      `@      W@      1@      .@      ;@     �F@       @      $@      9@      ,@      1@      5@      :@      D@       @              8@      Q@               @     �L@      &@     @U@     �H@     @Q@      F@      @              @      ;@              @      0@      �?     �I@      ,@      7@      .@                      5@     �D@              @     �D@      $@      A@     �A@      G@      =@      @      �?     @V@     �h@      "@      &@     �`@      4@     ��@      >@     �z@     �^@      @      �?      N@     �`@              �?      V@      &@     P}@      1@     �r@     @T@      �?              &@     �D@                      .@       @     �g@      @     @R@      *@                       @      =@                      $@       @      _@      @     �K@      (@                      @      (@                      @             �P@              2@      �?              �?     �H@      W@              �?     @R@      "@     `q@      ,@     @l@      Q@      �?      �?      H@     �U@              �?      M@      "@      n@      *@      h@     �P@      �?              �?      @                      .@              C@      �?     �@@       @                      =@     @P@      "@      $@     �F@      "@      d@      *@     �_@     �D@      @              7@      P@      "@      @     �F@      @      d@      *@     @_@     �D@      @              1@     �J@      @      @     �A@      @     �`@      &@     �U@      :@       @              @      &@      @       @      $@              ;@       @      C@      .@      �?              @      �?              @               @                       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��2z-@�	           ��@       	                   �5@7���@k           Z�@                           �?bG�֞�@�           ��@                           �?�|��@�           ؆@������������������������       ��\��WE@�            �q@������������������������       �:ވ/�v@           �{@                           �?�Nd-!@�            0v@������������������������       �_g9��@U             a@������������������������       �$ZF�)@�            `k@
                           �?���AT	@�           ��@                          �:@���(��@           �|@������������������������       �[��I@�            �r@������������������������       ��֌G@^            �c@                          �7@Ȯ�Dtr	@�            �@������������������������       ���t�`�@�            �h@������������������������       ��i�m(�	@0           �}@                          �7@֝����@2           p�@                           @Ŏ��j@6           @�@                           �?Y�}yL@G           ��@������������������������       �X�����@3           �~@������������������������       ��s�*E�@           �z@                          �3@��*�:�@�            �w@������������������������       ��W�$g@�            �i@������������������������       �l�b�@k            �e@                           @�XAk��@�            �x@                            �?$j���&@K             [@������������������������       ��T}��@+             M@������������������������       �h�|��@              I@                           @a !�h@�             r@������������������������       �W����@(             Q@������������������������       �t��+@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@     Ȃ@      >@     �F@     �z@     �W@     p�@     �j@     ��@     Pv@      9@      3@     �i@     �w@      2@     �B@     pr@     @R@     `y@     �e@     �u@     �n@      6@      @     �S@     �f@       @      0@     @`@      9@     p@      Q@     �i@     @Y@      @      @     �M@      ^@      @      &@     �Z@      4@     `c@     �B@     �`@      R@      @      �?      "@     �J@       @      @      E@      @     �R@      1@     �L@      3@              @      I@     �P@       @      @      P@      .@      T@      4@     @S@     �J@      @              3@     �O@      @      @      8@      @     �Y@      ?@     @R@      =@                      $@      7@      @       @      (@      �?      C@      3@      1@      &@                      "@      D@      �?      @      (@      @      P@      (@      L@      2@              (@     �_@     �h@      $@      5@     �d@      H@     �b@     �Z@     �a@     �a@      0@      @     �E@     �S@      @      @     �P@      2@     �L@      >@     �P@     @S@      @             �A@      J@      @      @      E@      @     �F@      6@      E@      G@      @      @       @      ;@              @      9@      ,@      (@       @      9@      ?@               @      U@     �]@      @      ,@     �X@      >@      W@      S@     @R@     �P@      $@      @      B@      F@              @      4@      @      7@      0@      <@      1@              @      H@     �R@      @      @     �S@      ;@     @Q@      N@     �F@     �H@      $@      �?     @T@     �k@      (@       @     �`@      6@     0�@      D@     �y@     @\@      @              M@     @f@      &@      @      T@      *@     �@      9@      s@     @R@      @              D@     �_@      @      @     �G@      @     �y@      1@      j@     �G@                      ;@     �H@              @      @@      @      n@      $@     �X@      8@                      *@     �S@      @              .@       @     �e@      @     �[@      7@                      2@     �I@      @      @     �@@      @     @`@       @      X@      :@      @              ,@      *@      @      @      *@              S@      @     �P@      &@      �?              @      C@      @              4@      @      K@      �?      >@      .@       @      �?      7@      E@      �?       @      K@      "@     @Y@      .@      [@      D@              �?      *@      "@                      2@       @      5@      �?      @@      &@                      @      @                      "@       @      (@              .@      $@              �?      @      @                      "@              "@      �?      1@      �?                      $@     �@@      �?       @      B@      @      T@      ,@      S@      =@                      �?      @              �?      *@       @      3@      @      0@      @                      "@      >@      �?      �?      7@      @     �N@       @      N@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJBK�LhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�y�?�j@�	           ��@       	                   �4@<�Ɲ=�@�           ��@                           @��H��@*           ��@                            �?y�:�[@V           ��@������������������������       ��
��'@)           0~@������������������������       ���`m��@-            �S@                           �?w��Z @�           ��@������������������������       �Tccz�?�            pq@������������������������       � ��_��@)           �}@
                           �?�=ƣ�Q@�           ��@                            �?d
�@.@           py@������������������������       �8�U�@�            �s@������������������������       �t����@:            @W@                          �<@J ���@�           P�@������������������������       �Ɍ����@<           (�@������������������������       ��k���@\            �a@                           �?�5K�7i@�           �@                           @��1��1@�            @u@                          �5@;l�E��@�            `n@������������������������       ��>d{�;@Y            `a@������������������������       ��0��%N@A             Z@                          �5@�3婕�?A            @X@������������������������       ���!.�?-            �O@������������������������       �`d6�<��?             A@                          �<@o�[�?	@           8�@                           @J.�A�	@�           h�@������������������������       ��/�`.�	@a           0�@������������������������       �Z��'�@h            �d@                           �?$G�f��@8            �V@������������������������       ��IE�@@             ,@������������������������       �
ۗc�@0             S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@      r@     ��@      =@      L@      |@     �T@     ��@     pp@     ȇ@     �w@      <@      @     �g@      x@      .@     �A@     0t@      I@     0�@     `g@     ��@     `o@      1@             �N@     @e@      @      $@     @]@       @     �}@     �R@     r@      Y@      @              >@     �T@               @      S@      @     �`@     �L@     �Z@     @Q@      @              =@     �R@               @     �N@              ^@     �H@     �U@     �L@      @              �?       @                      .@      @      (@       @      4@      (@                      ?@     �U@      @       @     �D@      @     �u@      2@     �f@      ?@                      @      7@               @      &@             �d@      @     �N@      @                      <@      P@      @      @      >@      @     `f@      (@     �^@      8@              @     @`@      k@      &@      9@     �i@      E@     �p@      \@     0q@     �b@      *@              <@     �M@      �?      @      G@      @     �[@      .@     �X@      A@      @              1@      G@      �?      @      ?@      @     @V@      $@     �R@      >@      @              &@      *@                      .@              5@      @      8@      @              @     �Y@     �c@      $@      6@      d@      B@     `c@     @X@      f@     @]@      @      @     �U@     @a@      "@      2@     �`@      ;@     �a@     �U@     �d@      U@      @              .@      3@      �?      @      ;@      "@      (@      $@      $@     �@@      @       @     �X@     @g@      ,@      5@     �_@     �@@      o@      S@     �h@     �_@      &@              8@      I@       @      @      B@       @     �]@      ,@     �N@      =@                      6@     �E@       @      @      A@       @      O@      ,@      B@      9@                      $@      6@              �?      4@       @      H@      @      2@      &@                      (@      5@       @       @      ,@              ,@      @      2@      ,@                       @      @              �?       @              L@              9@      @                      �?      @              �?                      C@              0@      @                      �?      @                       @              2@              "@                       @     �R@      a@      (@      1@     �V@      ?@     ``@      O@      a@     @X@      &@      @      L@     @]@      (@      ,@      T@      =@      `@     �J@      `@     @U@      &@      @     �H@     �X@      (@      ,@      Q@      8@      S@     �G@      T@     �Q@       @              @      3@                      (@      @      J@      @      H@      .@      @      @      3@      3@              @      &@       @      @      "@       @      (@                      �?                       @       @       @                       @      @              @      2@      3@              �?      "@              @      "@      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ#�2shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @X�<1@�	           ��@       	                    �?N�!.��@�           f�@                            �?x�*��z@�           �@                          �8@�u'�T@�            �h@������������������������       �燎���@b             b@������������������������       ��c�*�@             K@                          �<@��5Y�@&           �{@������������������������       ����@            x@������������������������       �-�V$�@$            �M@
                          �3@cn���:	@�           Ę@                           @���1��@           p{@������������������������       �&�n��#@�             i@������������������������       �#��?�J@�            �m@                           @��2�aj	@�           �@������������������������       ��Ӱ7	@f           ��@������������������������       �̡�d�@g            �d@                          �4@�����@+           X�@                           �?�/Cm@A           ��@                            �?�Q�w��?�            �u@������������������������       �n?���?5             V@������������������������       �eK�d�?�             p@                           @�^��>m@g           ��@������������������������       ��[��tH@:            �W@������������������������       �E����@-           �}@                           @ާ/��@�            �@                           @{�v�@�           ��@������������������������       ��'�+r�@^           ��@������������������������       �U���-@�             h@������������������������       ����A�@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        $@     �r@      �@      >@     �E@     �|@     @U@     �@     `m@     ��@     �v@      @@      $@      k@     �t@      5@      C@     t@      P@     @w@     �h@      x@      o@      ;@      �?      L@     �S@              @     @R@      @      d@      D@      c@     �N@      @      �?      "@      ?@                      0@      @     �H@      @     �N@      4@      @               @      4@                      (@      @      E@      @     �H@      @      @      �?      �?      &@                      @              @      �?      (@      1@                     �G@     �G@              @     �L@      @      \@      A@      W@     �D@      @              C@     �D@              @     �H@      @      [@      <@     �U@      7@      @              "@      @               @       @              @      @      @      2@              "@      d@     @o@      5@     �@@      o@     �L@     `j@     �c@     �l@     �g@      4@       @     �@@      Q@      @      @      M@      @     �[@      A@      P@      I@      @              &@      B@      @      @      :@      �?     �F@      &@      A@      :@               @      6@      @@                      @@      @     @P@      7@      >@      8@      @      @      `@     �f@      1@      ;@     �g@      J@     @Y@     �^@     �d@     @a@      .@      @      \@     �b@      0@      6@     �c@      H@      W@      V@     �c@      ^@       @      @      0@      ?@      �?      @      ?@      @      "@      A@       @      2@      @              T@      k@      "@      @     `a@      5@     x�@     �C@     0y@     �\@      @              C@     �\@       @      �?      F@      @     �{@      ,@     �j@     �D@      �?              .@      A@                      (@             @j@      @     �P@      @      �?                      @                       @             �P@              (@       @                      .@      =@                      $@             �a@      @     �K@       @      �?              7@      T@       @      �?      @@      @      m@      &@     `b@     �B@                      $@      (@                      @       @      :@      @      7@      &@                      *@      Q@       @      �?      :@      �?     �i@      @      _@      :@                      E@     �Y@      @      @     �W@      2@     �j@      9@     �g@     @R@      @             �D@     �Y@      @      @     �V@      *@     �j@      7@     �g@     @R@      @              2@      U@      @      @     �L@      *@      e@      3@     �b@      H@                      7@      2@      �?      �?     �@@              F@      @     �C@      9@      @              �?              @              @      @      �?       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��j�j@�	           ��@       	                     �?^DE ��@           ܓ@                          �8@m����@�           ��@                          �3@]	�B�@Y           x�@������������������������       ��5���	@�            �q@������������������������       �˥�Z0@�            0q@                          �?@�đ��@S             `@������������������������       ��"$�/�@L            �]@������������������������       ����N�@             $@
                          �5@ɸ����@f           8�@                            @}Н�@�            �w@������������������������       �1D��ͨ�?a            @b@������������������������       �݌椧x@�             m@                          �7@�\���@�            �i@������������������������       �ǥ����@&             N@������������������������       �[i�h�@Z             b@                            @�D�8SU@�           ��@                          �5@ ���@�           x�@                           @�#X� x@�           ��@������������������������       ��s��@H           �@������������������������       ����!�@O            ``@                           @���v"	@           ��@������������������������       �P4ڙ�	@:            @������������������������       ���2E<@�            �t@                          �@@��EE� 	@�           ��@                           �?nC����@�           �@������������������������       ��@�#l@�            �r@������������������������       ���'a��@-           �{@������������������������       ���W�@	             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     `s@      �@      3@     �P@     �|@     �T@     ؎@     �m@      �@     Px@      ?@      �?      T@     �e@      @      0@     �]@      &@     |@     �D@     Pr@      U@      @      �?     �I@     �Z@      �?      $@     �J@      @     �k@      0@      d@      M@       @              G@     �S@      �?      @     �E@       @     `i@      *@     �`@      ?@                      3@      F@              �?      &@              ]@      @     �Q@      2@                      ;@      A@      �?      @      @@       @     �U@      "@      P@      *@              �?      @      =@              @      $@      @      2@      @      :@      ;@       @      �?      @      <@                       @      @      2@       @      :@      :@       @               @      �?              @       @                      �?              �?                      =@     @P@       @      @     @P@      @     �l@      9@     �`@      :@      �?              1@      <@              @      A@       @      g@      *@     �S@      0@      �?              @       @                      .@              V@      @      8@       @      �?              *@      4@              @      3@       @     @X@      "@     �K@      ,@                      (@     �B@       @       @      ?@       @     �E@      (@     �J@      $@                      "@      $@                      @      �?      &@              4@      @                      @      ;@       @       @      9@      �?      @@      (@     �@@      @              0@     �l@     �u@      0@     �I@     @u@     �Q@     Ѐ@     �h@     �@     s@      <@      &@      d@     �n@      @      =@     �l@     �I@     �y@     �b@     �v@     �j@      0@      @     �O@     �c@      @      (@     @\@      ,@     @r@     �P@      l@     �Y@      @       @     �I@     `a@      @      &@     @Y@      @     p@      L@     �j@     �T@      @      @      (@      1@              �?      (@      $@     �A@      &@      $@      4@              @     @X@      V@      @      1@     @]@     �B@     �^@     @T@     `a@     �[@      (@      @      N@     �J@       @      .@     �Q@      >@     �E@      N@      S@     @R@      $@             �B@     �A@      �?       @     �G@      @     �S@      5@     �O@      C@       @      @     �Q@      Y@      $@      6@     �[@      4@      _@      H@     �a@      W@      (@      @     @Q@      Y@       @      6@     �[@      4@      _@     �E@     �a@     �U@      (@       @      ?@     �C@      @      &@      F@      @     �D@      @     �N@      G@      @      �?      C@     �N@      @      &@     �P@      .@     �T@      B@      T@     �D@      @       @      �?               @                                      @       @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���[hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?+�� �D@�	           ��@       	                     �?<��]Y@           �@                           @��@&��@�            Pu@                          �;@�~zj@�            `k@������������������������       ���wB��@�            @j@������������������������       ��ӿ� @             "@                           �?�]�I��?H            �^@������������������������       �Bۖ1M��?!            �L@������������������������       ���Uݭ� @'            @P@
                           �?�'�U��@C           8�@                          �<@��DY��@:           �~@������������������������       ��98�@'           �|@������������������������       ���2h�.@             ;@                          �<@�$�!��@	           �{@������������������������       ��!8S��@�            y@������������������������       ��7�g�@             F@                          �6@��4l B@�           ��@                           @L�L��+@           x�@                           @[��J� @           ��@������������������������       �t���v�@�           ��@������������������������       ����Q@S           ��@                           �?&<��^@             ?@������������������������       �k{��0J@             *@������������������������       �G\�s��@
             2@                           @��I��Y	@�           x�@                            �?��'���	@�           ��@������������������������       �I0A@�`
@�            �m@������������������������       ����@�^	@           `z@                          �<@aWշ�@�            �u@������������������������       �� s���@�            `r@������������������������       �<4)��@#             K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �p@     ��@      :@      M@     �~@     @W@     ��@     `j@     X�@     @v@      <@             �S@      g@      @       @     @]@      $@     �|@     �@@     �q@     @X@      @              &@      J@      �?       @      9@      @     `a@      @     @T@      4@      �?              &@      C@               @      5@      �?     �O@      @      N@      1@      �?              $@     �B@               @      2@             �O@      @      N@      ,@      �?              �?      �?                      @      �?                              @                              ,@      �?              @       @      S@      �?      5@      @                               @                                     �E@              &@      �?                              (@      �?              @       @     �@@      �?      $@       @                     �P@     �`@       @      @      W@      @     t@      ;@      i@     @S@      @              ?@      Q@       @      @     �H@      @      g@      2@     @W@     �A@                      >@     �O@       @      �?     �G@      @     �f@      1@     @V@      :@                      �?      @              @       @               @      �?      @      "@                      B@      P@               @     �E@       @      a@      "@      [@      E@      @              ?@     �M@                     �@@       @     �`@      @     @Z@      >@      @              @      @               @      $@              @      @      @      (@              1@     �g@     @x@      7@      I@     �w@     �T@     8�@     @f@     @     0p@      8@      &@     �Z@     �m@      @      6@     @h@     �C@      z@     �X@     pu@     �a@      &@       @     @Z@     �m@      @      6@     �g@     �@@      z@      X@     0u@     �`@      &@      @     @P@     @c@       @      *@      a@      :@     �p@     �G@     �n@      Y@      @      �?      D@     �T@      @      "@      K@      @     �b@     �H@     @W@     �A@      @      @      �?       @                      @      @       @       @      @       @              @      �?                               @      @      �?      �?               @                               @                      �?      @      �?      �?      @      @              @      U@     �b@      1@      <@     �f@      F@     �`@      T@     @c@      ]@      *@      @     �O@     @Z@      .@      6@     @_@     �D@     �J@     �P@     �Q@      T@      *@              4@      ?@      @      .@     �B@      3@      5@     �@@      9@      8@      @      @     �E@     �R@      $@      @      V@      6@      @@     �@@     �F@      L@      @              5@      F@       @      @      M@      @      T@      ,@      U@      B@                      .@     �C@              @      C@      @     @S@      ,@     @S@      9@                      @      @       @              4@              @              @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?~E�f�[@�	           ��@       	                    �?��2<ٸ@�           �@                           �?���@�           ��@                          �8@��I�0�@�            @m@������������������������       �Ƭ;: �@o            �e@������������������������       �!���~�@&             O@                            �?����ku @            {@������������������������       �@\)	��?C            �X@������������������������       ���z��� @�            �t@
                           @G��c�@c           H�@                          �7@Xf3:�@�            0u@������������������������       �Raˈl@�            �m@������������������������       �\�(V�*@=             Y@                          �2@�JL�4@�            �j@������������������������       �I9����?=            �V@������������������������       �hg��T@P             _@                          �4@��1W6@�           �@                           �?TU��@�           ��@                          �1@��]��-	@           @z@������������������������       �r#o�;@C             [@������������������������       ���~x�	@�            �s@                          �1@ܲ�A@�            �@������������������������       ��v��x�@�            pp@������������������������       ��u��q�@:           �@                            �? ���@�           p�@                           @2��U/	@�           ��@������������������������       �\k�ڤ	@<           @�@������������������������       ��dQOɪ@�            �p@                           @�Az�L�@�           P�@������������������������       ���#F"	@+           �|@������������������������       �@Ji3K@�            �o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �s@     Ѐ@      9@      K@     �|@     �V@     ��@      m@     `�@      v@     �B@      �?      S@     `c@      @      &@      [@      &@     �{@      D@     pq@     �T@       @      �?     �C@     �R@      @      &@      N@      @     Pq@      3@     �`@      D@              �?      8@     �@@      @       @      @@      �?      I@      0@      C@      ;@                      ,@      ;@      @       @      4@      �?     �G@      (@      =@      0@              �?      $@      @              @      (@              @      @      "@      &@                      .@      E@              @      <@      @     `l@      @     @X@      *@                              @                      @      @     �L@              6@       @                      .@     �B@              @      8@      @     @e@      @     �R@      @                     �B@      T@      �?              H@      @     �d@      5@      b@     �E@       @              ?@      I@                      B@      �?      R@      2@     �W@      >@      @              ;@     �@@                      6@             �J@       @     �R@      6@                      @      1@                      ,@      �?      3@      $@      4@       @      @              @      >@      �?              (@      @     �W@      @      I@      *@      �?              @      @                      �?              K@       @      3@      @      �?               @      9@      �?              &@      @     �D@      �?      ?@      "@              (@     �m@     �w@      4@     �E@     �u@     �S@      �@      h@     P@     �p@      =@      @     �T@     �d@      @      0@      ^@      ,@     �u@     �Q@     �n@     �[@      &@      @      D@     �H@      @      @     �Q@       @     �O@      B@      P@      O@      &@      �?      @      3@      �?      �?      .@              8@      @      3@      3@              @      A@      >@      @      @     �K@       @     �C@     �@@     �F@     �E@      &@              E@      ]@      �?      "@      I@      @     �q@     �A@     �f@      H@                       @     �C@              �?      (@             �\@      (@     �O@      *@                      A@     @S@      �?       @      C@      @     @e@      7@     @]@     �A@              @     �c@     @k@      .@      ;@     �l@     @P@     �l@     �^@     p@     �c@      2@      @     �U@     @[@      @      2@     �]@     �D@     @\@     �T@     @_@      S@      &@      @     �M@      R@      @      .@      U@      B@      G@     �Q@     �Q@     �I@      $@              ;@     �B@      �?      @      A@      @     �P@      &@     �K@      9@      �?      @     �Q@     @[@      &@      "@     �[@      8@     �\@      D@     �`@     �T@      @      @      M@      T@      "@      @     @R@      6@     �F@     �B@     @P@      N@      @              *@      =@       @      @     �B@       @     �Q@      @     �P@      7@      @�t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��SwhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @y�'�gA@�	           ��@       	                   �:@`ѫ���@Y           �@                           �?�~"�NW@a           �@                           �?`̘t��@\           p�@������������������������       �$�l�c�@�            �o@������������������������       ���R6��@�             s@                           @����M	@           T�@������������������������       ���w���@�           4�@������������������������       �߂����@Y             a@
                           @��(�6V	@�            �x@                          �<@-m��Q	@�             r@������������������������       ��|6��	@G            �]@������������������������       ��g���@n             e@                          �=@|����@C             [@������������������������       �8Ӕ�}�@&             M@������������������������       �Jf�>@             I@                            @��$G@<           �@                            �?XF�f�p@�           L�@                           �?Dl��|@�             v@������������������������       �
���7��?H            @Z@������������������������       � �\��@�             o@                           @c��)��@�           Đ@������������������������       �Gj�~A@�            �@������������������������       �1��.�@�            �p@                           @3�pu0V@�            pr@                          �4@�;]� @�            `l@������������������������       �Jё&2@I            @`@������������������������       �4�n�G�?9            @X@                           @`$�R�@*             Q@������������������������       ��\8��?             7@������������������������       �]���W@            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     Ps@     ؁@      <@      D@     �{@      W@     Ў@     �j@     ��@     @v@     �@@      0@     �k@     pt@      4@      <@     �r@      R@     �v@     �e@     0x@     �n@      >@      @      f@     �q@      .@      9@     p@     �L@     �t@     �`@     pt@     @d@      6@              K@     @T@       @      @     �R@      @      c@      9@     ``@      =@      �?              4@     �D@       @      @     �E@      @     �Q@      1@      C@      *@      �?              A@      D@                      @@      �?     �T@       @     @W@      0@              @     �^@     �i@      *@      6@     �f@      J@     `f@     �Z@     �h@     �`@      5@      @     @[@      g@      *@      6@      c@     �C@      d@     @W@     �g@     @^@      *@      �?      *@      5@                      >@      *@      2@      ,@      @      (@       @      &@      G@     �D@      @      @      G@      .@      B@      D@      N@     @U@       @      @      B@     �C@      @      �?     �E@      "@      4@      3@      I@      J@      @      @      ,@      .@      @              1@      @      (@      @      =@      $@      @              6@      8@      �?      �?      :@      @       @      ,@      5@      E@      @      @      $@       @               @      @      @      0@      5@      $@     �@@      �?      @      @                      �?       @              (@      "@      @      7@                      @       @              �?      �?      @      @      (@      @      $@      �?      �?     �U@     �n@       @      (@      b@      4@     X�@     �D@      {@     @[@      @      �?     �R@     �l@      @      (@     @^@      3@      @     �C@      u@      W@      @              3@     �I@                      9@      @      d@      "@     �P@      4@                              .@                       @       @     �P@              1@      @                      3@      B@                      7@       @     �W@      "@     �H@      1@              �?     �K@      f@      @      (@      X@      .@      u@      >@     �p@      R@      @      �?      C@     �]@              @      R@      "@     �q@      4@      i@      I@       @              1@     �M@      @      @      8@      @      J@      $@     @Q@      6@      �?              *@      0@      @              7@      �?     @^@       @     �X@      1@                      "@      ,@                      ,@              X@       @     @T@      &@                       @      (@                      $@             �J@       @     �D@      @                      �?       @                      @             �E@              D@      @                      @       @      @              "@      �?      9@              1@      @                      @                              @              (@                      �?                               @      @              @      �?      *@              1@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��K�I@�	           ��@       	                   �1@i	��@a           .�@                           �?NN���@�           ��@                           �?њ0.��@t            �g@������������������������       ��L7�@5             U@������������������������       ����X��@?            �Z@                            @u�J�� @           P{@������������������������       �C!S�@�            0v@������������������������       ���#��X�?/            �T@
                           �?E�@�           ��@                          �3@|2@G           X�@������������������������       ���K��@�            r@������������������������       �����@�            @m@                            @�+���i@�           d�@������������������������       �XM���@�           ��@������������������������       �Y�G�q@�            0r@                          �<@��B-�@O           Ț@                           �?7�5'c�@{           l�@                            �?����T@�            `v@������������������������       �,�{��[@y            �h@������������������������       ���w�@j            @d@                           �?��^�u@�           ��@������������������������       ��rj�@           �y@������������������������       �M(ڈ�$@�           Ȃ@                          @A@�� D	@�            pu@                           @�<�?@�@�            �s@������������������������       �$�l'�@�            �o@������������������������       �Eu���@)            @P@                           �?�e�b��@             8@������������������������       �B8iY�o @             (@������������������������       �_�z|�X@             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     0�@      ;@     �K@     �~@     @S@     �@     �k@     @�@     �u@      B@      "@     @Z@     `s@      ,@      ;@     �o@      :@     �@     �X@     �~@      b@      1@              1@     �T@      �?      @     �L@             p@      :@     �a@     �C@       @              "@      ?@      �?       @     �C@              E@      *@      A@      3@                       @      (@                      4@              =@      @      *@      @                      @      3@      �?       @      3@              *@       @      5@      0@                       @      J@               @      2@             �j@      *@     �Z@      4@       @              @      E@               @      2@             �d@      @     �V@      4@       @              �?      $@                                      H@      @      1@                      "@      V@     `l@      *@      7@     �h@      :@     |@     @R@     �u@     @Z@      .@             �B@     @R@      �?      @     �C@      @     `h@      2@     �]@      ?@                      6@      A@               @      (@      @     �\@      @      S@      5@                      .@     �C@      �?      @      ;@      �?     @T@      *@      E@      $@              "@     �I@     @c@      (@      0@     �c@      6@     �o@     �K@     �l@     �R@      .@      �?      D@     �]@      @      (@     �Y@      (@     @h@      E@     @e@     �I@      "@       @      &@     �A@      @      @      L@      $@      N@      *@     �M@      7@      @       @     �f@      n@      *@      <@      n@     �I@     r@     �^@      t@     @i@      3@       @      b@     �g@      &@      2@     �h@     �@@     `p@     �U@     �q@     �_@      .@              ?@      G@      �?      �?     �C@      @     @Z@      .@     @W@      3@      @              .@      8@                      9@              O@      @      I@      $@      @              0@      6@      �?      �?      ,@      @     �E@       @     �E@      "@               @     �\@     �a@      $@      1@     �c@      <@     �c@     �Q@     @h@     �Z@      (@      �?      D@     �K@      @       @     �O@       @     �M@      ;@     �T@     �K@      &@      �?     �R@     �U@      @      "@      X@      4@     �X@      F@      \@      J@      �?      @     �A@      J@       @      $@     �E@      2@      ;@     �B@     �@@      S@      @       @      <@     �H@       @      $@     �C@      0@      ;@      B@     �@@     @R@      @       @      5@      A@       @      "@      ;@      ,@      .@      B@      9@     @P@      @              @      .@              �?      (@       @      (@               @       @              @      @      @                      @       @              �?              @                      @       @                      @                      �?              �?              @       @      �?                      �?       @                               @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJӽ�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�y��qN@�	           ��@       	                    �?���X�o@           ؒ@                          �8@�{UN�@�           ��@                            �?�n�Gk@F           �@������������������������       ��AJk�� @Q             _@������������������������       ��AZ�U�@�            Px@                           �?�@fsY@Q            �]@������������������������       �f	�T�@-            �P@������������������������       �K�yjp@$            �I@
                          �<@��|���@y           ��@                          �2@G� �@W           0�@������������������������       �t�i��Y @�            �h@������������������������       �v���͆@�            �s@                          �?@Ö�7PO@"            �L@������������������������       ������~@             C@������������������������       ��.q�;�?             3@                          �:@���U�8@�           &�@                           �?$I�˖�@�           ܡ@                            @,���@c             e@������������������������       ��5�D��@@            �Z@������������������������       �b7WA�@#             O@                           @�P��,c@R           ��@������������������������       �i>Y���@�           ��@������������������������       �@JDZh@@a           0�@                           �?A�2�z	@           Pz@                            �?9�+���	@�            @n@������������������������       ���I��@*            �P@������������������������       ���<S�	@j            �e@                           @X*؃�@p            `f@������������������������       ��w��D	@             G@������������������������       ����u�@S            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     �@      <@     �K@     �{@     �T@     �@     �l@     �@     0v@      <@      �?     �S@     �c@      @      (@     �[@      &@     �z@      C@     0r@      R@       @      �?     �E@     �Q@       @       @     �O@       @     �m@      6@      a@      E@                      A@     �M@       @      @     �J@      @     @j@      ,@     �\@      2@                               @              @      3@      �?      L@       @      @@      @                      A@     �I@       @      @      A@       @     @c@      (@     �T@      .@              �?      "@      &@               @      $@      @      :@       @      6@      8@              �?       @      @               @      $@      �?       @      @      &@      0@                      �?      @                              @      2@      @      &@       @                     �A@     @V@      �?      @     �G@      @      h@      0@     `c@      >@       @              >@     @U@      �?      �?     �@@      @     @g@      $@     �b@      3@      �?              @      6@              �?      "@             �Y@      @      G@       @                      7@     �O@      �?              8@      @      U@      @     �Y@      &@      �?              @      @              @      ,@              @      @      @      &@      �?              @      @                      @              @      @      @      "@      �?              �?      �?              @      &@              �?                       @              5@     �k@     0x@      9@     �E@     �t@     �Q@     ��@     �g@      �@     �q@      :@      "@     �f@     pu@      0@      ?@     p@     �L@     ��@      c@     `~@      i@      8@      @      2@      7@              &@      >@      @      0@      2@      ?@      .@               @      $@      "@              @      4@      �?      .@      @      ;@      $@              �?       @      ,@              @      $@       @      �?      &@      @      @              @     `d@      t@      0@      4@     `l@      K@     �@     �`@     p|@      g@      8@      @     �\@      i@      *@      &@     `c@     �G@     �j@     @\@     @g@      Z@      5@              H@     �]@      @      "@      R@      @     �r@      6@     �p@     @T@      @      (@      D@      F@      "@      (@     @R@      ,@      B@      C@      M@     �T@       @      (@      4@      ;@      "@       @     �A@      (@      ,@      6@      7@      M@       @      �?      �?      @              @      (@      @      @      $@      @      *@      �?      &@      3@      5@      "@      @      7@      @      @      (@      0@     �F@      �?              4@      1@              @      C@       @      6@      0@     �A@      9@                      �?       @              @       @      �?      @      @      @      $@                      3@      "@                      >@      �?      3@      "@      ?@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���8�G@�	           ��@       	                    �??����[@[           �@                          �4@�u�6S@�           `�@                            �?+X��$3@�           �@������������������������       �kz$&�)@�            `u@������������������������       ������@�            pr@                           �?�2��U)@F            �[@������������������������       ��)R�@(            �M@������������������������       ��P4G��@             J@
                           �?�ڋY�@�           $�@                           @%Ó	@E           �@������������������������       ��g�Ef�@;            @������������������������       �tT^Rv�@
             ,@                          �4@��]�z�@A           X�@������������������������       �u#�]O@�           Ї@������������������������       �j�!y�@^             b@                           �?�a����@L           P�@                           �?�gj�Ų	@           x�@                          �<@p�_���@�            `l@������������������������       �oV{�w�@n            �f@������������������������       �y~~�}�@              G@                           �?A�����	@}           `�@������������������������       ���\��	@|            `g@������������������������       ���c?�	@           y@                           @e�7@A           (�@                           @�����@�           ��@������������������������       �@�U@u           ��@������������������������       ��o��j@�             l@                            �?_	aK��@E             ]@������������������������       �<U%h�@"             N@������������������������       ��<��^�@#             L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     pr@     0�@      7@     �K@     @|@     @W@     �@     �l@     P�@     pv@      ?@      $@     @^@     0r@      @      7@     �j@      @@     ��@     �U@     @@     �b@       @              A@      [@              @      F@      @     �s@      0@      h@      @@      �?              =@     �S@              @      D@      @     �p@      ,@      e@      <@      �?              4@     �F@               @      >@             �`@      @     �W@      "@                      "@      A@               @      $@      @      a@      @     �R@      3@      �?              @      =@                      @       @     �D@       @      8@      @                       @      .@                       @       @      7@              (@      @                      @      ,@                       @              2@       @      (@      �?              $@     �U@     �f@      @      3@      e@      ;@     �y@     �Q@     @s@     �]@      @      $@     �K@      P@      @      &@      W@      2@     �T@      E@     @Q@      N@      @       @     �I@     �O@      @      &@     �V@      .@     �T@      E@     @Q@     �M@      �?       @      @      �?                      �?      @                              �?       @              @@     �]@      @       @      S@      "@     �t@      =@     �m@     �M@      @              <@      X@      @      @      M@      @     �r@      7@     `h@     �J@                      @      7@               @      2@      @     �@@      @      F@      @      @       @     �e@     `l@      1@      @@      n@     �N@     s@     �a@     `s@      j@      7@      @     @X@     @Y@      (@      3@     �a@      D@     �R@     �S@     �Z@     �^@      3@              ;@      @@      �?      @      F@      �?      @@      (@     �F@      7@      @              8@      7@      �?       @      D@      �?      <@      &@     �C@      "@      @              @      "@              @      @              @      �?      @      ,@              @     �Q@     @Q@      &@      (@      X@     �C@     �E@     �P@     �N@     �X@      0@       @      0@      9@       @      @      @@       @      7@      (@      3@     �A@      @      @      K@      F@      "@      @      P@      ?@      4@     �K@      E@      P@      $@      @     @S@     �_@      @      *@      Y@      5@     �l@      P@     �i@     �U@      @      @      N@     @Z@       @      *@     �U@      2@     @j@      E@     `h@     @T@       @      @      I@      R@               @      L@       @     �e@     �A@      _@     �M@       @              $@     �@@       @      @      >@      $@     �A@      @     �Q@      6@                      1@      5@      @              ,@      @      4@      6@      "@      @       @               @      @       @              @      @      $@      2@      @      @                      "@      0@      �?              &@              $@      @      @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ^K�.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�'T@�	           ��@       	                   �5@ ��?=	@
           �@                           �?�fH�@            �@                           �?���.@�            �q@������������������������       ���k]@@            �\@������������������������       �~���7@e            @e@                           @����@_            �@������������������������       �q��]#@�            �v@������������������������       �Da�%S�@r            �f@
                           �?�,�6��	@            �@                           @�Dq݊�@�             q@������������������������       ������@f            �c@������������������������       �U����@L            �\@                           �?���7�J
@T           ��@������������������������       ������
@�            �j@������������������������       ������A
@�            �u@                           �?ؕ�TC@�           ��@                            @������@�            �@                           @+k��j@l           ��@������������������������       �h���@X            �a@������������������������       �r_|
@            {@                           @�H�;�?Q            @`@������������������������       �E�	V�@             B@������������������������       ���k���?;            �W@                           @U�IR�@�           �@                          �7@�ڠC�@d           �@������������������������       ������@�            �@������������������������       �J�x��@�             v@                          �8@�I	�:/@{            `h@������������������������       �`�Q6�5@X             a@������������������������       �C��V�@#             M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     ��@      >@     �O@     �|@     �S@     ��@     `j@     ��@      v@      ;@      6@      f@     �m@      6@     �B@     �m@     �G@      p@     �`@     �q@      h@      4@      @     �S@      Y@      @      (@     �]@      1@     �f@     �I@     @d@     �W@      @              6@     �@@      �?      �?      =@      @     @U@      2@     @R@      3@                      @       @                      .@              B@      @      D@      @                      2@      9@      �?      �?      ,@      @     �H@      &@     �@@      .@              @     �L@     �P@      @      &@     @V@      ,@      X@     �@@     @V@      S@      @      @      C@      F@      @      @      N@      $@      L@      .@     @R@     �K@      �?       @      3@      7@       @      @      =@      @      D@      2@      0@      5@      @      0@     �X@     @a@      .@      9@     �]@      >@     �R@     �T@      _@     @X@      0@      @      <@     �D@       @      @      F@       @      E@      4@     �F@     �A@      @      @      1@      *@                      ;@              @@       @     �@@      6@      �?              &@      <@       @      @      1@       @      $@      (@      (@      *@       @      (@     �Q@     @X@      *@      3@     �R@      <@     �@@     �O@     �S@      O@      *@      @      6@     �G@      @      @      6@      &@      ,@      5@     �@@      7@      @      "@      H@      I@      @      *@     �J@      1@      3@      E@      G@     �C@      @             @^@     0t@       @      :@      l@      @@     ��@     @S@     �@     @d@      @              6@     @W@       @      @      G@      @     `t@      @      d@     �@@      @              3@     @V@       @      @      A@      @     �o@      @     �_@      =@      @              @       @               @      @      @      L@       @     �H@       @       @              ,@     @T@       @      �?      =@      @     �h@      @     @S@      5@      �?              @      @               @      (@             �Q@              A@      @                      �?       @                      "@              &@              $@      @                       @       @               @      @              N@              8@      �?                     �X@     �l@      @      5@     @f@      9@     �z@     �Q@     v@      `@      @              T@      i@      @      1@     �c@      5@     0x@      H@     �s@     �[@      �?             �G@     �c@      @      *@     �Z@      ,@     pt@      ;@     �l@      Q@      �?             �@@     �E@      �?      @      J@      @      N@      5@     �V@     �E@                      3@      >@      �?      @      4@      @     �C@      6@     �A@      2@      @              @      9@              @      $@       @     �A@      2@      3@      0@      @              ,@      @      �?              $@       @      @      @      0@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJcC�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@����P|@�	           ��@       	                    @�i�n�@^           *�@                           �?
5[{t@@
           |�@                          �4@._!�ZL@A           0�@������������������������       ���YD@�            Ps@������������������������       ��F���o@~             j@                           �?`J����@�           d�@������������������������       ��F|`�d	@�            �v@������������������������       ��t�^̓@�           X�@
                           �?�ޏ3L@T           ؔ@                           @��3��?+           }@������������������������       ��2�`���?�            �s@������������������������       �
>*���?[            �b@                           @ӎ4>��@)           (�@������������������������       ���ţ@u            �f@������������������������       �^'��@�           ��@                            @���(0S	@O           ��@                            �?�����@�           ��@                           @4Y�2T�@4           �~@������������������������       ��5ǔ�	@�            �t@������������������������       �zg��t�@b             d@                           �?������@Z            �a@������������������������       �4J���@            �G@������������������������       ��w�ν�@>            �W@                           �?R1�ʢ�	@�            �s@                           �?S�D}�	@�            �j@������������������������       ���ۄU;@9            �W@������������������������       �Q ᄯ	@I            �]@                          �=@�/^��@?             Z@������������������������       �Z�J9<�@2            @T@������������������������       �?\qC#@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �s@     �@     �@@     �E@     P}@      X@     X�@     �k@     ��@     `w@      =@      1@     @j@     �x@      4@      =@     @v@      M@     h�@     @`@     H�@     `n@      .@      0@     �b@      n@      1@      3@      o@      D@     �s@      [@      s@     @c@      .@             �A@     �P@      �?      @      M@      @     `d@      6@     �_@     �@@      @              ,@     �D@              @     �@@       @     @W@      5@     �R@      ;@      �?              5@      9@      �?      @      9@      @     �Q@      �?      J@      @       @      0@     @\@     �e@      0@      *@     �g@     �A@     �c@     �U@     �f@     @^@      (@      @      E@     @R@      "@      @     �L@      (@     �H@      >@      @@     �F@      @      $@     �Q@     �Y@      @      "@     �`@      7@     �Z@      L@     �b@      S@      @      �?      O@      c@      @      $@      [@      2@     p�@      6@     pu@     @V@                      (@      L@              �?      8@             �m@      @      [@      3@                      (@      B@                      3@              f@      @     �M@      &@                              4@              �?      @              O@      @     �H@       @              �?      I@      X@      @      "@      U@      2@     �q@      0@     `m@     �Q@              �?      0@      :@       @              ,@      (@      N@      @      B@      &@                      A@     �Q@      �?      "@     �Q@      @     `l@      *@     �h@     �M@              "@     @Z@     @^@      *@      ,@     @\@      C@     �_@      W@     �e@     ``@      ,@      @     �P@      S@       @      @     �U@      <@     �R@     @P@     �^@     �U@      &@      @      G@     �O@      �?      @     �L@      8@     �L@     �M@     �W@     �Q@      @      @      9@     �J@      �?      @      D@      7@      D@     �A@      K@     �G@      @       @      5@      $@               @      1@      �?      1@      8@      D@      7@      @              4@      *@      �?      �?      =@      @      2@      @      <@      1@      @              &@      @                      "@      �?      @               @      "@      @              "@       @      �?      �?      4@      @      (@      @      :@       @              @     �C@     �F@      &@       @      ;@      $@     �I@      ;@      I@      F@      @      @      >@      B@       @       @      6@      $@      .@      7@      =@     �@@      @       @      ,@      0@      @      �?      *@      @      �?       @      3@      0@       @      �?      0@      4@      @      �?      "@      @      ,@      5@      $@      1@      �?              "@      "@      @      @      @              B@      @      5@      &@                      "@      @      @      @      @              =@      @      1@      @                              @                                      @      �?      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��_zhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @E��h�;@�	           ��@       	                   �9@$�9�@m           V�@                           �?�nS�	@#           4�@                           �?ZRLFq@�           ��@������������������������       ��q�.�@5           ~@������������������������       ��f|�*	@�           0�@                           �?##�bb@6           `~@������������������������       ��Q)��@            �i@������������������������       ��}D�u�@�            �q@
                           �?��wN�	@J           ��@                          �<@����R@X            �b@������������������������       �	v^��@'             N@������������������������       ���ۙ�>@1            �V@                           �?�2Ov��	@�            �x@������������������������       �fq���`@;            @W@������������������������       ��9)�
@�            �r@                          �4@���!I@&           x�@                           @�54�@K           ؍@                           �?�� ��@�            �i@������������������������       ��S�4	�@F            �Z@������������������������       �'�;jQ @=            �X@                            �?����� @�           h�@������������������������       �Ҥ�L)�?]            �a@������������������������       ����q��@k           ��@                          �6@��L�"@�           �@                           @�F�}Ő@�            Pq@������������������������       �ࢯ��t@�            �o@������������������������       ���鴄@             8@                           @h���g@-           �|@������������������������       �MQ8f@           z@������������������������       ��"+��+@            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �p@     ��@      <@      N@      {@     �S@     x�@     `n@     X�@     w@      :@      .@     �g@     `u@      5@      G@     �r@     �L@     �w@      h@     x@     �p@      4@      @     @a@     �o@      *@     �A@     �j@      @@      u@     �`@     pt@     @f@      (@      @      [@     �g@      &@      8@     �d@      9@     �g@     �Y@     �k@     @a@      "@       @     �@@     @T@              @     �P@      @     �X@     �A@     @Z@     �G@       @      @     �R@      [@      &@      1@     �X@      5@      W@     �P@     �]@     �V@      @              >@     �P@       @      &@      G@      @     @b@      ?@      Z@      D@      @              &@     �@@       @      @      5@      @      N@      "@      C@      5@      @              3@     �@@              @      9@      @     �U@      6@     �P@      3@              "@     �J@     �U@       @      &@      U@      9@      G@      N@      M@     @W@       @      @      *@      8@              @      <@      �?      5@      2@      .@      6@       @      @      @      ,@                      &@      �?      (@      @      @                              @      $@              @      1@              "@      (@       @      6@       @      @      D@     �O@       @       @      L@      8@      9@      E@     �E@     �Q@      @              @      *@      �?              7@      @      "@      @      *@      6@      �?      @     �B@      I@      @       @     �@@      5@      0@     �B@      >@     �H@      @      �?     �S@     �l@      @      ,@     @a@      5@     ��@      I@     �z@     �X@      @             �A@     �[@      @      @     �G@      @     �{@      5@     �m@      G@                      &@      H@                      &@      @     @T@      @     �A@      "@                      "@      ;@                      @             �A@      @      .@       @                       @      5@                      @      @      G@              4@      �?                      8@      O@      @      @      B@             �v@      .@     @i@     �B@                      @      @              �?       @             @V@              <@      @                      4@     �K@      @      @      <@              q@      .@     �e@      @@              �?     �E@      ^@       @      @     �V@      0@     �f@      =@     �g@      J@      @               @     �J@      �?      �?      C@       @     @V@      �?     �L@      0@      @               @      I@      �?      �?     �@@      @      V@      �?     �J@      *@                              @                      @      @      �?              @      @      @      �?     �A@     �P@      �?      @     �J@       @     �W@      <@     �`@      B@      �?      �?      9@     @P@      �?      @      H@       @     �U@      4@     �^@     �A@                      $@       @                      @               @       @      $@      �?      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�B�YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�0�pt@�	           ��@       	                    �?����>	@�           ��@                           �?�Af�O\@2           @~@                           �?�����@|             i@������������������������       �y�I���@9            @V@������������������������       ��g���S@C             \@                            @`'�4�x@�            �q@������������������������       ���a1@j@^            �b@������������������������       ��8�3��@X            �`@
                           @�ni�	@�           ��@                           �?�"
�,o	@�           p�@������������������������       �۷�K:�@            y@������������������������       �{����	@�           `�@                             @���@            �A@������������������������       ����%��?             8@������������������������       ��� 8��@             &@                          �7@��g��@�           L�@                          �4@D`����@H           ��@                          �1@!���@�           �@������������������������       �+ۀ�@           �z@������������������������       �؄8%�@�           h�@                          �5@(��v� @Q           p�@������������������������       �	����@�            `m@������������������������       ��W#�c@�            0t@                          �<@ʭt���@q           ��@                           �?�$�*x@$           �|@������������������������       ��u~�>@�            `k@������������������������       �"Q�!��@�             n@                           @�C^	�a@M            �\@������������������������       �n���h@.            �P@������������������������       ���m�@             H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pq@     @�@      B@     �E@      |@     @S@     0�@     `i@     ��@     u@      @@      1@     �c@     �m@      5@      ;@     @o@     �C@     �n@     @\@     �o@     �f@      ;@             �E@     �Q@       @       @     �P@      �?      \@      6@     @Z@     �J@      �?              1@      <@                      5@             �L@      @      M@      1@                       @      &@                      &@              7@      @      6@      &@                      "@      1@                      $@              A@              B@      @                      :@      E@       @       @      G@      �?     �K@      3@     �G@      B@      �?              .@      3@                      9@      �?      ;@      $@     �@@      4@      �?              &@      7@       @       @      5@              <@      "@      ,@      0@              1@      ]@      e@      3@      3@     �f@      C@     �`@     �V@     `b@      `@      :@      *@     �[@     �d@      3@      3@     �f@     �A@     �`@      U@      b@      `@      1@       @      9@     @R@       @      "@     @Q@      *@     �O@      8@      P@      L@              &@     @U@     �W@      1@      $@     @\@      6@     @Q@      N@     @T@     @R@      1@      @      @       @                      �?      @      �?      @       @              "@      �?      @                              �?                      @                      "@      @               @                              @      �?               @                      �?     �]@     �s@      .@      0@      i@      C@     ��@     �V@     ��@     `c@      @              S@     @o@      *@      &@     �_@      8@     8�@     �G@     �{@     �X@       @             �H@     �d@      @      @     �R@      @     @@     �A@     �r@     �Q@                      ,@      K@              @      3@              i@      $@     �Z@      4@                     �A@      \@      @      @      L@      @     �r@      9@     �g@     �I@                      ;@      U@      @      @     �I@      5@     `f@      (@     �a@      <@       @              @      >@               @      5@      *@     �Q@      @     �S@      @       @              5@      K@      @       @      >@       @      [@      @     @P@      5@              �?      E@     �O@       @      @     �R@      ,@      \@     �E@      d@      L@      @      �?      :@      G@       @      @      M@      (@     �X@     �A@      a@     �C@       @      �?      (@      5@               @      >@             �F@      0@     �R@      0@       @              ,@      9@       @       @      <@      (@      K@      3@      O@      7@                      0@      1@              �?      0@       @      *@       @      8@      1@      �?               @       @              �?      (@       @       @       @      &@      ,@      �?              ,@      "@                      @              @              *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJI�GGhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�.mMb@�	           ��@       	                    �?����I	@�           |�@                           �?t��JDm@1           0~@                           �?_4����@q            �f@������������������������       �W@��@2            @S@������������������������       ���C�E@?             Z@                            @օ�0E@�            �r@������������������������       �D"G%��@f            `d@������������������������       �O���@Z            `a@
                          �:@�gx��	@�           �@                           @mef�\	@4           ��@������������������������       ��C+�@`           0�@������������������������       �S�j���	@�            `u@                          �?@m$]�i�	@�             l@������������������������       ��m��	@w            �f@������������������������       �h�B@�@             E@                           �?����J�@�           ԡ@                          �=@%�)D�@�           ��@                            @ ��n@�           L�@������������������������       �fh�]��@H           ��@������������������������       �?8oj+@{            `h@                           @@�4��ɧ@             =@������������������������       �����~��?             ,@������������������������       ��XV���@             .@                           @�C�=�@�           �@                            �?K�JY�@�            0u@������������������������       �(-A��@G             ]@������������������������       �n���@�            �k@                           @.Ȓ�3@�           8�@������������������������       �׿&9�@�           H�@������������������������       �d���@7            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     @r@      �@      C@     �G@     P{@     @V@     �@     �n@     X�@     @w@      ;@      .@     `e@      m@      >@      ;@     �n@      H@     @j@     �b@     @q@      i@      7@             �G@     �T@      @      @     �O@      @     @W@      =@     @X@      J@      @              *@      >@                      2@             �J@      @      D@      4@       @              @      "@                      @              ;@      @      3@      "@                      "@      5@                      (@              :@       @      5@      &@       @              A@      J@      @      @     �F@      @      D@      8@     �L@      @@      @              2@      9@               @      ?@      @      1@      "@     �B@      .@      @              0@      ;@      @      @      ,@      �?      7@      .@      4@      1@              .@      _@     �b@      ;@      6@     �f@      E@     @]@     �^@     `f@     �b@      1@       @      Z@     �`@      0@      4@      c@      >@     @Z@     �V@     @c@      Y@      (@       @     �J@     �R@      &@      *@      Y@      4@     @P@      F@      ^@      S@      @      @     �I@     �L@      @      @      J@      $@      D@     �G@      A@      8@      "@      @      4@      3@      &@       @      ?@      (@      (@      ?@      9@     �H@      @      @      0@      ,@      @              8@      (@      (@      :@      3@     �D@      @      �?      @      @      @       @      @                      @      @       @              �?     @^@     ps@       @      4@     �g@     �D@     x�@      X@     ��@     `e@      @      �?      K@     �c@      @      *@     @[@      2@     y@      A@     �o@     @W@      �?      �?     �G@     @c@      @      *@     @Z@      *@     y@      ?@     @o@      V@      �?      �?      G@     �`@       @      (@     @V@       @     �t@      <@     �h@      P@      �?              �?      5@      �?      �?      0@      @      R@      @     �I@      8@                      @      @                      @      @              @       @      @                      @                              @                      @              @                      @      @                              @                       @       @                     �P@     @c@      @      @     �T@      7@     �w@      O@     �q@     �S@      @              ;@     �H@              @      ?@      "@     �T@      ;@     @T@      ;@       @              @      .@               @      @      @      @@      $@      8@      ,@       @              6@      A@              �?      :@       @     �I@      1@     �L@      *@                      D@     @Z@      @      @     �I@      ,@     �r@     �A@     @i@     �I@      �?              =@     �V@      @      @      G@      *@     �q@      9@      g@      C@      �?              &@      .@       @              @      �?      3@      $@      2@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ڪVhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?OiZ�@�	           ��@       	                    �?�}U�@           ��@                          �;@H+���T@)           ~@                            �?&��_n@           `z@������������������������       �mo0�n�@U             b@������������������������       ���$��7@�            `q@                           �?B��&@#            �M@������������������������       ���u�2@            �@@������������������������       �:;�?�@             :@
                            �?d�"�U	@�           p�@                          �4@��/�\�@�            �u@������������������������       �#�X���@K            @]@������������������������       �w���^	@�            �l@                           �?S�%��O	@            �@������������������������       �E)4�G@�            pt@������������������������       ��w9�(�	@<           �@                          �4@r�R@�@�           ��@                           �?1�9=w�@�           �@                            @_��� @           �z@������������������������       ��J��[6@�            �u@������������������������       ��s&��?1            �S@                          �1@ �y�?�@�           Ј@������������������������       �B
dc^o@�            p@������������������������       ����+�@G           Ȁ@                           @d��s@�           $�@                          �5@ϔ����@�           x�@������������������������       �����R@P             ]@������������������������       �WK���{@D           �@                            �?1��[@           �y@������������������������       �bc@=            @T@������������������������       ���H �@�            �t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      s@     P�@      ;@     �J@     �}@      S@     (�@     �i@     ��@     `t@      4@      1@      e@     `r@      0@     �A@      p@      G@     @n@     �`@     �p@      e@      .@       @      G@      X@      �?      $@      L@       @      ^@      1@     @V@     �D@      �?             �B@      V@      �?      @      I@       @     �\@      .@      U@      8@      �?               @     �E@                      *@              C@      @     �@@      @                      =@     �F@      �?      @     �B@       @     @S@      &@     �I@      3@      �?       @      "@       @              @      @              @       @      @      1@               @      �?      @              @       @              @       @      @      (@                       @      @               @      @               @               @      @              .@     �^@     �h@      .@      9@      i@      F@     �^@     �]@     @f@      `@      ,@       @     �E@     �E@      @      (@      M@       @      B@     �H@     �N@      >@      @              1@      @                      .@      �?      2@      .@      <@      ,@       @       @      :@      B@      @      (@     �E@      @      2@      A@     �@@      0@      �?      *@      T@     `c@      (@      *@     �a@      B@     �U@     @Q@     @]@     �X@      &@      �?      9@     @Q@       @      @     �K@       @      E@      9@     �D@      H@      @      (@     �K@     �U@      $@      @     �U@      <@      F@      F@      S@      I@      @             �`@     @r@      &@      2@     �k@      >@     ��@      R@     X�@     �c@      @             �H@     @c@      @      $@     �X@      @      @      >@     �r@     �Q@      �?              ,@      I@              @      9@             �j@      @     �W@      3@      �?              (@      G@               @      7@             �e@      @      P@      2@      �?               @      @              �?       @             �B@              ?@      �?                     �A@      Z@      @      @     �R@      @     �q@      8@     �i@      J@                      @      ?@              @      .@             �\@      @      Q@      0@                      =@     @R@      @      @     �M@      @     @e@      4@     @a@      B@                     �U@     @a@       @       @     �^@      9@     0p@      E@     �o@     �U@      @             �P@     �Q@      �?      @     �T@      4@     @d@      >@     �`@      G@      @              @      2@                      1@      @      8@      @      ?@      @      @             �M@     �J@      �?      @     �P@      *@     @a@      ;@     �Y@     �D@                      4@     �P@      @       @      D@      @     @X@      (@      ^@      D@                      @       @       @              $@      �?      6@      @      2@      $@                      1@     �M@      @       @      >@      @     �R@      @     �Y@      >@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��mMhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@LTFE7F@�	           ��@       	                    �?�WN4Ȅ@X           �@                           @-�SE�@�           �@                           �?�@���@�            �t@������������������������       �ti��]O@X            @a@������������������������       ����N��@}            `h@                           �?�;C���@	            y@������������������������       �Z�z^o@s            �e@������������������������       �N���y�@�            @l@
                           �?�c�t�@z           ��@                           �?y;�\�@�           Ȇ@������������������������       �I�]^�?�            �q@������������������������       �c����@            |@                           �?x��U�@�           p�@������������������������       ���,��� @�            `m@������������������������       ��.�溴@'           0~@                           @�BϪ'�@Q           �@                          �;@�Z���p	@�           L�@                           �?�)z� �@�           �@������������������������       ��S�갢@�             i@������������������������       ��6"?uo	@v           ��@                          �>@t��9_�	@�            `s@������������������������       ��9�L��@�            @i@������������������������       �x�=5
	@G             [@                           �?�F�P"@�           ��@                          �9@D&0Mn�@�             s@������������������������       �rE4O{@�            `h@������������������������       �1�!�@A            @[@                          �<@��z,@�             t@������������������������       �J��@�            �o@������������������������       �{@HKÕ@%             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `t@     ��@      ;@     �O@     @{@      R@     ��@     �k@     ��@     �v@      7@      @      `@     Ps@      @      9@      k@      ?@     8�@     �V@     P�@      d@      @      @      L@      [@      @      &@     �X@      .@      b@     �K@     @c@     �S@      @      @      @@     �F@              �?      @@      �?     �U@      9@     �T@      9@      �?      �?      @      (@                      *@             �D@      $@     �G@      &@               @      =@     �@@              �?      3@      �?     �F@      .@     �A@      ,@      �?       @      8@     �O@      @      $@     �P@      ,@     �M@      >@      R@     �J@      @              &@      :@              @      3@      @     �B@      &@     �@@      9@               @      *@     �B@      @      @     �G@       @      6@      3@     �C@      <@      @              R@      i@      @      ,@     �]@      0@     ��@     �A@      w@     �T@       @              ;@     �W@              @     �T@      @     �q@      1@     �d@     �G@      �?              *@      ;@              @      6@             `d@       @     �E@      @                      ,@     �P@              �?     �N@      @      ^@      .@     @^@     �D@      �?             �F@     �Z@      @       @      B@      "@     `o@      2@     �i@     �A@      �?              $@     �@@                      "@              \@       @     �L@      @      �?             �A@     �R@      @       @      ;@      "@     `a@      $@     `b@      >@              *@     �h@     �o@      4@      C@     `k@     �D@     �r@     @`@     �r@     `i@      0@      *@     @c@      f@      0@      :@     �c@     �@@     @^@     @Z@     @c@      a@      ,@      @     �]@      `@      (@      3@     �]@      4@     @Z@     @R@     �]@      R@       @              B@     �@@      �?      �?      9@       @     �I@      @     �B@      @      �?      @     �T@     �W@      &@      2@     @W@      2@      K@     �P@     �T@     �P@      @      "@     �A@     �H@      @      @      D@      *@      0@      @@     �A@      P@      @      @      4@     �C@      @      @      5@      (@      (@      "@      6@     �J@       @      @      .@      $@      �?      @      3@      �?      @      7@      *@      &@      @              F@      S@      @      (@     �N@       @     �f@      9@     @b@     �P@       @              <@      H@              "@      7@       @     �V@      "@      R@      5@       @              0@      A@              @      1@       @     �I@       @     �G@      5@       @              (@      ,@              @      @             �C@      @      9@                              0@      <@      @      @      C@      @     �V@      0@     �R@      G@                      *@      7@       @       @      4@      @     �T@      ,@      Q@      7@                      @      @       @      �?      2@               @       @      @      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�؉MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����B6@�	           ��@       	                    �?��o��@�           l�@                          �<@��=��@�           `�@                           �?(��^�V@z           �@������������������������       �Ac�3G6@	           py@������������������������       ����g�@q            `e@                            �?���c�v@-            �R@������������������������       �-��a� @             4@������������������������       ����o�@"             K@
                          �3@U
Mi�6	@�           ��@                           @�Uo�5�@           @|@������������������������       �d�@f&�@�             m@������������������������       �޼cw	<@�            `k@                           �?�Ā��	@�           ��@������������������������       ���
�@�            �p@������������������������       �BȾQ�r	@           Њ@                          �7@��^�%�@.           L�@                           �?�jY�@           ��@                            �?4³iޜ @8           �}@������������������������       ��3�: @�            @p@������������������������       ����L�K @�            `k@                           @�4�8��@�           8�@������������������������       �ξ؈)?@           @z@������������������������       ��\S�9@�            0v@                           @��ㅢ�@           �z@                           @(��FeL@B             [@������������������������       �ѷ���@#             L@������������������������       ��?��2m@             J@                           @j͗��@�            t@������������������������       �]�o�.%@0            �R@������������������������       �*��@@�            �n@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     `r@     ��@      =@     �H@     @{@     �T@     �@      m@     �@     �u@     �A@      *@     �l@     @u@      8@      A@     `r@     �O@     �x@     �g@     px@     �l@      ?@      �?     �O@     �S@       @      "@     �R@       @      d@     �@@     �b@     �P@      @      �?     �L@     �P@       @      @     �P@       @     @c@      :@     �a@      G@      @      �?      E@     �L@       @      @      K@      @      V@      :@      W@      ?@      @              .@      "@              �?      *@      @     �P@             �H@      .@                      @      (@              @      @              @      @      "@      4@       @               @       @                                                      @      @       @              @      @              @      @              @      @      @      .@              (@     �d@     `p@      6@      9@     �k@     �K@      m@     �c@      n@     @d@      8@       @      6@     �P@              @      O@      @     �]@     �G@     �S@     �C@      @      �?      *@      C@              @     �@@             �O@      (@     �G@      4@              �?      "@      <@              �?      =@      @     �K@     �A@      @@      3@      @      $@     �a@     �h@      6@      2@     �c@      J@     �\@     �[@     @d@     �^@      1@              *@      G@      @       @      B@      &@      E@      4@     �F@      C@      @      $@     @`@     �b@      2@      $@     �^@     �D@     @R@     �V@     @]@     @U@      (@      �?     �P@      l@      @      .@     �a@      3@     ؃@     �E@     �y@     @]@      @             �G@     @e@      @      $@     @V@      1@     ��@      2@     �r@     @Q@       @              0@      L@      �?       @      :@       @     `o@      @     @Y@      0@       @              @      E@      �?              *@       @     ``@      �?      K@      &@                      &@      ,@               @      *@              ^@      @     �G@      @       @              ?@     �\@      @       @     �O@      .@     pq@      (@     �h@     �J@                      2@      I@       @              =@       @     �d@      $@      [@      >@                      *@      P@      �?       @      A@      @     �\@       @     @V@      7@              �?      3@     �K@      �?      @     �J@       @     @Z@      9@     @\@      H@       @      �?       @      .@              �?      7@              8@      �?      :@      .@              �?       @      ,@                      @              *@              $@      $@                              �?              �?      1@              &@      �?      0@      @                      1@      D@      �?      @      >@       @     @T@      8@     �U@     �@@       @              @      @                      @      �?      3@      "@      .@      ,@       @              &@      B@      �?      @      :@      �?      O@      .@      R@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJb��GhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @a����/@�	           ��@       	                    �?��
wK�@�           R�@                           �?���87@�           ��@                          �1@���
>�@2           �}@������������������������       �t��v��@2            �S@������������������������       ������*@            �x@                            �?�ýr�@u             h@������������������������       ���}���?*             O@������������������������       �#7e;�&@K            @`@
                           �?f6��A	@�           D�@                           �?!�q.'@G             [@������������������������       ��$8	�@             =@������������������������       �3Yg��@3            �S@                            �?Ť�w$	@�           ��@������������������������       �� �<��@           �{@������������������������       �kK�Bx-	@�           0�@                            @�Z1�=@7           ��@                          �4@��=9�p@�           D�@                           @Tp��5@�           h�@������������������������       ��m磭� @           8�@������������������������       ��S�s�@q            �d@                           @����5@�            �@������������������������       � �m�:�@�           ��@������������������������       �����@
             0@                           �?���5�@�            �p@                           @.,AU�?I            @\@������������������������       �B��?             A@������������������������       ��e�]d�?4            �S@                          �6@�e�~@`            �c@������������������������       �de��� @;            @W@������������������������       �ߥI,9@%            @P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     ��@      =@     �J@     �|@     @T@     h�@     �h@     x�@     �v@      =@      ,@     `i@     �v@      :@     �B@     �s@     �K@     x@     �d@     pw@     �o@      8@      �?      P@     �Y@      �?      @     �T@      @      e@      >@     �`@     @Q@      @      �?     �H@     �T@      �?      @     �O@       @      X@      9@     �V@      K@      @              @      "@                      &@             �@@      @      *@      @              �?      G@     �R@      �?      @      J@       @     �O@      4@     @S@      I@      @              .@      4@                      3@      �?      R@      @     �F@      .@                       @      $@                      �?      �?      ;@              3@       @                      *@      $@                      2@             �F@      @      :@      *@              *@     `a@     p@      9@      @@     �m@      J@      k@     �`@      n@      g@      5@       @      .@      .@              $@      7@      @       @      $@      0@      (@                      @      &@                      @       @               @       @       @               @      $@      @              $@      2@      �?       @       @      ,@      $@              &@      _@     @n@      9@      6@     �j@     �H@     �j@     @_@      l@     �e@      5@      �?      A@     @R@      @      @     @Q@      "@      U@      H@     @P@      D@      *@      $@     �V@      e@      5@      .@      b@      D@     ``@     @S@     �c@     �`@       @             �W@     �n@      @      0@      a@      :@     `�@      A@     �y@     �Z@      @              V@     `k@      @      ,@     @[@      9@     �@      ?@     �t@     �V@      @             �C@     �Y@      �?      @     �B@             �u@      0@     @g@     �G@       @              =@     @S@               @      4@             Pr@      $@     �b@      B@                      $@      9@      �?      @      1@             �I@      @      C@      &@       @             �H@     @]@       @      @      R@      9@     �d@      .@      b@      F@      @             �G@     @]@              @     @Q@      3@     �d@      *@      b@      F@      @               @               @              @      @      �?       @                                      @      ;@               @      <@      �?     �[@      @     �S@      .@                      @      (@              �?      @              L@      @     �@@       @                      �?      $@                                      *@              $@                               @       @              �?      @             �E@      @      7@       @                      @      .@              �?      9@      �?      K@             �F@      *@                      @       @                      ,@      �?      A@              @@      �?                      �?      @              �?      &@              4@              *@      (@        �t�bub�       hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJip@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @I &Wd@�	           ��@       	                    �?���9�@c           �@                          �;@#��z�[@�            �@                            �?'�2���@{           ��@������������������������       �� ��@�@~             i@������������������������       �O��Mn@�            �x@                           �?^�[�>@2            �T@������������������������       ��2�6=@(            �Q@������������������������       �m�:.1�@
             *@
                          �2@�(Kb^�	@�           t�@                            @ViR��@�            �r@������������������������       �G��Yq@k            �e@������������������������       �@�:�Ex@I            �_@                           @�����	@           Ē@������������������������       ���0^��	@�           Ȉ@������������������������       ��ꁔh�@           �y@                           @�dB##@?            �@                            �?����N@�           l�@                          �1@E'�2D@�           0�@������������������������       ���T��?c            �c@������������������������       ����ٱQ@0           �~@                          �<@N3s���@Q           ��@������������������������       �n���g@>           @������������������������       ��@b��@             B@                            �?(RoG�[@[           h�@                          �5@��h�r�@I             `@������������������������       �3��c�l�?#            �O@������������������������       ����^@&            @P@                          �6@��G�:@           �z@������������������������       �����@�            �q@������������������������       �f���Q@\             b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     8�@      =@     �L@     �z@      V@     ��@     �k@     @�@     `y@      ?@      .@     @i@     �s@      2@      G@     �r@     �P@     `v@     �f@     w@     Pq@      =@       @     @Q@     �Y@      �?      @     �R@      @      d@      5@      c@     �S@      @              N@     @W@      �?      @     �O@      @     @c@      1@     @a@     �K@      @              &@     �B@              �?      8@      �?      H@      @     �M@      ,@      �?             �H@      L@      �?      @     �C@      @     �Z@      (@     �S@     �D@       @       @      "@      "@               @      &@              @      @      ,@      8@       @       @      @       @               @      $@              @      @      &@      7@                       @      �?                      �?               @      �?      @      �?       @      *@     �`@     �j@      1@      D@      l@      O@     �h@     �c@      k@     �h@      8@      �?      8@      C@              @     �E@      @      Q@      ?@     �I@      @@      @      �?      1@      8@                      5@      @      E@      9@      7@      *@      @              @      ,@              @      6@       @      :@      @      <@      3@              (@     @[@      f@      1@     �B@     �f@      L@     @`@      `@     �d@     �d@      5@      "@      T@     @\@      0@      7@     �]@     �G@     �R@     �O@     �^@      \@      ,@      @      =@      P@      �?      ,@     �O@      "@      L@     @P@     �E@      K@      @             �W@     @m@      &@      &@     �`@      5@     x�@      D@     p{@      `@       @             �P@     �b@      �?      @      R@      1@      }@      <@     pr@     @S@      �?              D@     �U@      �?              ;@      (@     `n@      ,@     �d@     �K@                      @      (@                       @             �T@              E@      *@                      B@     �R@      �?              9@      (@      d@      ,@     @_@      E@                      ;@     �O@              @     �F@      @     �k@      ,@      `@      6@      �?              9@     �O@               @      ?@      @     �j@      (@      _@      4@      �?               @                      @      ,@              "@       @      @       @                      ;@      U@      $@      @      N@      @     �c@      (@      b@      J@      �?              "@       @      @      �?      $@       @     �F@      @      A@      &@                              @              �?      @             �A@              0@      @                      "@      @      @              @       @      $@      @      2@      @                      2@      S@      @      @      I@       @      \@       @     �[@     �D@      �?              @      L@      @       @      <@       @     �U@       @     �R@      4@      �?              &@      4@      �?      @      6@              9@      @     �A@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�pHhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�"��k@�	           ��@       	                    �?�4���@t           8�@                           �?�m�X��@�           ��@                          �<@ ���@k             f@������������������������       ��g���@a             d@������������������������       �+�%W�@
             0@                          �<@�P�!�@6           0~@������������������������       �ܦ7k��@           �z@������������������������       ������@#            �J@
                          �4@����A�	@�            �@                           �?����@p           0�@������������������������       �(���p�@�            �w@������������������������       �,ޙ^u@y             i@                          �:@` @��	@c           �@������������������������       ���SE�	@�           ��@������������������������       ���5�`	@�            �t@                           �?%	J�<@C           ��@                            �?*��+T@q           ��@                          �6@�#����?S            @`@������������������������       ���ۇ�?@             Y@������������������������       ���l�t@             >@                           @�j���~@            {@������������������������       �+|�@@�            �l@������������������������       ��0��Y@�            �i@                          �8@����L@�           �@                           �?kD�d@8           ��@������������������������       �h�we	m@$            �K@������������������������       ����@           ��@                            �? B��@�             m@������������������������       �@�T�&@"             I@������������������������       �32�Pz�@x            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     ��@     �D@     �F@     �}@     @T@     ��@     �l@     ��@     �w@      ;@      1@     �h@     �t@      >@     �@@      u@     �P@     �v@      h@     �v@     �n@      9@              H@     �T@       @      @     @V@      @     `f@      A@     �c@      K@      @              $@      5@                      8@             �K@      @     �K@       @      �?              @      2@                      6@             �J@      @     �K@      @      �?              @      @                       @               @                      @                      C@      O@       @      @     @P@      @      _@      ?@     @Y@      G@       @             �B@     �M@       @      @     �J@      @     �^@      6@     @X@      <@                      �?      @               @      (@               @      "@      @      2@       @      1@     �b@     �n@      <@      :@     �n@      O@     `g@     �c@      j@      h@      6@      @     �D@     �T@      @      $@     @W@      (@     �Z@     �M@     @W@     @Q@      @      @      A@      C@      @       @     �Q@       @     �K@      B@     �N@     �N@      @              @      F@      �?       @      6@      @     �I@      7@      @@       @              (@      [@     �d@      6@      0@     @c@      I@     @T@     �X@      ]@      _@      0@      @      U@     �]@      *@      *@      Z@     �@@      K@     �M@     �S@      K@      *@       @      8@     �F@      "@      @      I@      1@      ;@      D@     �B@     �Q@      @       @      X@     �m@      &@      (@      a@      ,@     �@      C@     Pz@     ``@       @              0@      U@      @              >@      @     �o@      @     @a@      9@                              @      @              $@      �?      R@              >@      @                              @                      @             �P@              4@      @                              @      @              @      �?      @              $@       @                      0@     @S@                      4@      @     �f@      @      [@      2@                      (@     �B@                      &@      @     �Z@      @      I@      @                      @      D@                      "@             @S@      @      M@      (@               @      T@      c@       @      (@     �Z@      $@     0v@      ?@     �q@     �Z@       @       @      J@     @`@      @       @     �R@      $@     t@      1@     �l@     @P@       @       @      @      &@                      @       @      *@      @      *@                             �H@     �]@      @       @     �Q@       @     @s@      $@     �j@     @P@       @              <@      6@      @      @      ?@              A@      ,@     �K@     �D@                       @      @                      @              &@      @      .@      $@                      :@      2@      @      @      <@              7@      "@      D@      ?@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�I�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�ǿ[@�	           ��@       	                    �?\1
_�@E           ��@                           @�"�Q�@�           Ȇ@                           �??Y����@�            �t@������������������������       �oۥR��@`            �c@������������������������       �����@t            �e@                          �4@Kz��t��?�            �x@������������������������       ��y<W`��?�             u@������������������������       �ഡ ��?              M@
                           @��{�6�@}           ��@                            �?�\�9�k@�           P�@������������������������       ���G�5=@�            `i@������������������������       ��Q��h�@?           �@                           @����@�           ؆@������������������������       �������@l             f@������������������������       �0��'�@M           X�@                           �?���G �@B           ,�@                           �??~�v�
@(           ȋ@                            �?�(�(@�            @r@������������������������       �)�)D@8            @V@������������������������       �_���ڋ@|            `i@                          �@@C�Mg/a
@t           ��@������������������������       �aə�4
@h           �@������������������������       ���}��9@             4@                           @ۃo��@           ��@                           @�ꎢ�@m            �@������������������������       ��|r�u@�            �x@������������������������       ��.�}c`@o            �f@                           @,m�J@�             q@������������������������       �7[�z�|@j             e@������������������������       ��L��C_@C            @Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        @@     Ps@     ��@      ;@     �D@     �|@     @S@     Ў@     �l@     ؉@     pv@     �@@      "@     @_@     �r@      &@      .@     `i@      :@     ��@     �Z@      �@      d@      .@             �C@     @X@       @      @     �C@       @     s@      9@     �e@      E@      @              <@     �E@       @       @      ;@       @     �Y@      4@      S@      >@      �?               @      7@       @      �?      0@       @      L@      .@      5@      *@      �?              4@      4@              �?      &@              G@      @     �K@      1@                      &@      K@              �?      (@             `i@      @      X@      (@       @              &@      E@              �?      @             �e@      @     @U@      (@       @                      (@                      @              >@              &@                      "@     �U@     �i@      "@      (@     �d@      8@     x@     �T@     @u@     �]@      (@      "@      K@     �Y@      @      @     �Z@      ,@     ``@      Q@     �`@      R@      $@              0@      >@                      <@      @      D@      .@     �E@      5@      @      "@      C@     @R@      @      @     �S@      $@     �V@     �J@     �V@     �I@      @              @@     @Y@      @      @     �L@      $@     �o@      ,@     �i@      G@       @              $@      @@                      .@      "@      P@      "@      >@      @                      6@     @Q@      @      @      E@      �?     �g@      @      f@     �C@       @      7@      g@     @m@      0@      :@     �o@     �I@     �r@     �^@     �s@     �h@      2@      5@     @[@     @_@      *@      5@      a@     �@@     �Y@      T@     @]@     �\@      1@       @      1@     �F@      �?      @      J@      @      I@      2@      E@      H@      @              @      (@              @      .@      �?      .@      @      1@       @       @       @      &@     �@@      �?      �?     �B@      @     �A@      &@      9@      D@      @      3@      W@      T@      (@      ,@      U@      <@      J@      O@     �R@     �P@      (@      *@     �V@     �S@      (@      *@     @T@      :@      J@      O@     �R@      O@      (@      @      �?       @              �?      @       @                              @               @     �R@     @[@      @      @     �]@      2@     @h@     �E@     �h@      U@      �?       @      A@     �Q@      �?       @      T@      1@     �c@      9@     �`@     �I@               @      ;@      F@                     �M@      &@     �`@      (@     �S@      <@                      @      ;@      �?       @      5@      @      :@      *@      L@      7@                     �D@      C@       @      @      C@      �?      B@      2@     �O@     �@@      �?              8@      1@              @      5@              6@      @      I@      ;@                      1@      5@       @              1@      �?      ,@      *@      *@      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�~	#hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�m|��m@�	           ��@       	                    �?z���d�@           X�@                          �;@IJ"���@�           ��@                           �?Y�!���@o           ��@������������������������       ��  ��@x            �g@������������������������       �(vy�E@�            Pw@                          �>@V�I� �@'             Q@������������������������       �l�;Y�l@             G@������������������������       ����z�@             6@
                          �<@�X��I\@|           ��@                          �2@+�=��@b           ��@������������������������       �����AC@�             j@������������������������       �b-@�             v@                          �>@n:�@             F@������������������������       ��.�b�@             7@������������������������       ��O�Nʄ�?             5@                            @d`|p$F@�           �@                           @��;��@�           |�@                          �:@E����k	@P           ��@������������������������       �Fʩk�	@�           І@������������������������       ��)�\2@w            @g@                           �? Q��G@k           X�@������������������������       ���}$�@)             M@������������������������       ���\���@B           ��@                           @M\��@�           ��@                           �?Y�TK�Z	@�           0�@������������������������       ��bw�M�@+            @R@������������������������       ���C�0	@W           �@                           @�>9�O]@m            �e@������������������������       ���1&m@d            �c@������������������������       ����d@	             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     0r@     ȁ@      =@      M@      {@     @V@     ��@     `m@     ��@     pw@      @@      �?     �U@     `e@      @      $@     @\@      (@     �{@     �B@     pq@     �R@       @      �?     �C@      S@      @       @     �F@      "@     �o@      :@     @^@      F@      @             �B@      O@      @      @      D@      @      o@      5@      [@      =@      @              4@      8@      @              0@      �?     �J@      0@      C@      ,@      @              1@      C@              @      8@      @     `h@      @     �Q@      .@              �?       @      ,@              @      @      @      @      @      *@      .@              �?              ,@              @      @       @       @              &@      "@                       @                               @      �?      @      @       @      @                     �G@     �W@      �?       @      Q@      @     @g@      &@     �c@      >@      @             �E@     @V@      �?       @      J@      @     `f@      @     �c@      :@      @              @      9@               @      3@             �V@      @      I@       @       @              B@      P@      �?             �@@      @      V@      @     �Z@      2@       @              @      @                      0@              @      @       @      @      �?              @      @                       @              @      @      �?      @      �?              �?       @                      ,@              @              �?                      2@     �i@     �x@      6@      H@     �s@     @S@      �@     �h@     P~@     �r@      8@      $@     �b@     �p@      &@      @@     @j@      K@     P|@     �`@     �u@     �i@      .@       @     �U@      a@      @      6@     @_@      E@     �a@     �Y@     �[@     �^@      (@      @     �R@     �^@      @      1@     �W@      9@     �`@     �S@      W@     �Q@      "@       @      (@      ,@      �?      @      >@      1@      @      8@      2@     �J@      @       @     �N@     �`@      @      $@     @U@      (@     �s@      @@     `m@     �T@      @       @      @      &@               @      �?      @      "@       @      1@      @                      L@     @^@      @       @      U@      "@     �r@      >@     @k@     @S@      @       @     �L@      `@      &@      0@     @[@      7@     �_@      P@     �a@     �W@      "@       @      J@     �[@      @      .@     @W@      7@     �R@      O@     @V@     @R@      @      �?      @      (@              @      (@      �?      @      4@      @      "@      �?      @     �G@     �X@      @      $@     @T@      6@      R@      E@     @U@      P@      @              @      3@      @      �?      0@              J@       @     �I@      6@       @              @      2@       @      �?      *@             �I@       @      G@      6@                      �?      �?       @              @              �?              @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ'��fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���� @�	           ��@       	                    �?�P��\�@           h�@                            �?z���@3           �@                          �;@�RRk@�            �p@������������������������       ������@�             l@������������������������       ���H@             F@                           �?֘��u@�            �m@������������������������       ������5@=            @\@������������������������       �.Y\��c@N             _@
                          �;@�ԪS�q	@�           ��@                           �?k���@W           ��@������������������������       ��?��@�            �w@������������������������       ��`�16Y	@c           ��@                            �?�!�oS?
@�            �i@������������������������       �X?D(zQ@&             P@������������������������       ����e�	@_            �a@                           �? L�ۺ�@�           ޡ@                          �4@�/�"�@�           8�@                           �? o��{�?            �|@������������������������       ���ω�7 @�            �n@������������������������       ��[i����?�            �j@                            @�?�'m@�            �s@������������������������       ����De�@�            `p@������������������������       ���#KU?�?"             J@                           @$���&@�           ��@                          �2@sM �7�@           �y@������������������������       ��n/q$@=             U@������������������������       �bG�P
@�            �t@                           �?�%��')@�           $�@������������������������       �a��}@M           8�@������������������������       ��E���@q           �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     Ѐ@      ,@     �N@     `}@     �S@     �@     �j@     8�@     �v@      >@      2@      c@     �n@       @      >@     0p@     �G@     @m@     `a@     �p@      i@      7@      �?      I@      V@       @      @      O@       @     �Y@      =@     @Z@     �L@       @      �?      <@      I@      �?      @      3@             �G@      .@      Q@     �A@       @              8@     �C@      �?      @      1@             �F@      *@      P@      1@       @      �?      @      &@                       @               @       @      @      2@                      6@      C@      �?       @     �E@       @      L@      ,@     �B@      6@                      @      2@      �?       @      .@       @      =@      @      8@      *@                      3@      4@                      <@              ;@       @      *@      "@              1@     �Y@     �c@      @      9@     �h@     �F@     ``@     �[@     `d@     �a@      5@      $@     �T@     @`@      @      1@     �e@      <@     �]@      U@     �b@     �Y@      0@              5@      O@      �?      "@      S@      @     �Q@      A@     �L@      E@      @      $@     �N@      Q@      @       @     @X@      5@     �H@      I@     �V@      N@      (@      @      5@      =@       @       @      8@      1@      (@      :@      .@     �D@      @              �?      (@              �?       @      @      $@      @      @      &@      @      @      4@      1@       @      @      0@      &@       @      3@      &@      >@      �?      �?     �a@     0r@      @      ?@     `j@      @@     Ȉ@     @R@     ؀@     `d@      @              @@     �W@      �?      @     �H@      "@     �v@      @      g@      >@       @              1@      D@              @      4@             �n@       @      \@      5@                      "@      5@              @      0@             `a@       @      E@      *@                       @      3@                      @             @Z@             �Q@       @                      .@      K@      �?              =@      "@     �]@      @      R@      "@       @              *@      K@      �?              9@      "@      W@      @     �K@       @       @               @                              @              ;@      �?      1@      �?              �?      [@     �h@      @      :@     @d@      7@     �z@     �P@     0v@     �`@      @             �@@     �Q@      �?      $@     �M@      (@     �T@      C@     �Q@     �B@      �?              �?      .@                      &@              ?@      .@      @      @                      @@     �K@      �?      $@      H@      (@      J@      7@     �P@      ?@      �?      �?     �R@     �_@      @      0@     �Y@      &@     �u@      =@     �q@      X@      @      �?      B@     �O@      �?      *@     �L@       @      c@      &@     @`@     �H@      @             �C@      P@      @      @      G@      "@     @h@      2@     @c@     �G@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�qpshG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?R���76@�	           ��@       	                    �?�k�2��@�           ��@                          �4@�]�{@~           P�@                           @a[��@�            �p@������������������������       �wA1=@|             i@������������������������       ���$�!@%            @Q@                           �?�AU0@�            �u@������������������������       �Sd6�|@@             [@������������������������       ��Q�`Q�@�             n@
                            �?o�-3z�	@�           �@                           @��}t(�	@:           �~@������������������������       �١[/I�	@�            �v@������������������������       ������@T             `@                           �?�']��@G           ��@������������������������       �c�N
�W@Y             c@������������������������       ��.L�[	@�            �w@                           @���@�           ��@                           �?P/��p�@t           ��@                            �? �����@k            `c@������������������������       ��Œ܉ @=             W@������������������������       �ڳ�\�V@.            �O@                          �4@���7�c@	           0x@������������������������       �ĕ3Y�R@}             h@������������������������       ���@�@�            @h@                          �5@L.lCC@9           �@                           �?0�m&�I@�           �@������������������������       � Z�2\�?�            �x@������������������������       �����tb@�           h�@                           �?+h#��@�           �@������������������������       �t��M�g@�            �s@������������������������       �y�����@�            `t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      r@     `�@      :@      L@     �|@     �Q@     p�@     �m@     Ї@     Px@      <@      1@      d@     �o@      1@      ?@     Pp@     �C@      p@     �a@      m@      k@      6@      �?     �@@     �X@      �?      .@     �X@       @      b@     �C@     �Z@      Q@      @      �?      (@      E@              �?      F@      �?     @S@      *@     �L@      6@              �?      @      9@                      @@             �O@      @      K@      2@                       @      1@              �?      (@      �?      ,@      "@      @      @                      5@     �L@      �?      ,@      K@      @      Q@      :@      I@      G@      @              @      1@                      *@             �@@      @      9@      $@      �?              1@      D@      �?      ,@     �D@      @     �A@      5@      9@      B@      @      0@     �_@      c@      0@      0@     `d@      ?@     @\@     �Y@     @_@     �b@      2@      @      P@     �M@       @      &@     �R@      2@     �L@     �P@      L@      N@      *@       @      F@     �H@      @      $@      J@      1@     �E@     �B@     �J@     �D@      "@      @      4@      $@      �?      �?      7@      �?      ,@      >@      @      3@      @      &@     �O@     �W@       @      @      V@      *@      L@      B@     @Q@      V@      @              1@     �A@      �?      �?      9@              8@      $@      .@      9@              &@      G@     �M@      @      @     �O@      *@      @@      :@      K@     �O@      @      �?     @`@      q@      "@      9@      i@      ?@     Ј@     �W@     ��@     �e@      @             �H@     �R@      �?      @     @P@      (@     @b@      D@     @Z@      F@      �?              2@      &@              �?      &@       @     @P@      @     �B@      @                      &@      @              �?      �?       @      F@       @      9@      �?                      @      @                      $@              5@      @      (@      @                      ?@     �O@      �?      @      K@      $@     @T@     �A@      Q@     �C@      �?              @      @@      �?       @      8@      �?     �M@      .@      A@      5@                      ;@      ?@               @      >@      "@      6@      4@      A@      2@      �?      �?     @T@     �h@       @      4@      a@      3@     @�@      K@     �z@      `@      @              E@     �_@      @      (@     �P@      @     �}@      6@     q@      I@      @              .@      F@              �?      0@      �?     �k@      @     @S@      .@       @              ;@     �T@      @      &@      I@      @     p@      3@     �h@     �A@      �?      �?     �C@      R@      @       @     �Q@      ,@      e@      @@      c@     �S@       @      �?      :@      D@              @      =@      �?      X@       @     �P@      F@       @              *@      @@      @      @     �D@      *@     @R@      8@     @U@     �A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ubhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@q���;E@�	           ��@       	                    �?�NֶҲ@^           &�@                          �1@˧E�u>@�           ��@                           �?���[@v            �h@������������������������       �g{��@6             W@������������������������       �a�)�@@            �Z@                          �4@���@m           ��@������������������������       �c�5�"�@           P|@������������������������       �~�|#�@Z            `b@
                           @ۖ��C@{           ԕ@                           @t�s��@�           (�@������������������������       �)f�� @@�            �t@������������������������       ���`�+@�            `q@                           @XY�:P@�           ��@������������������������       �`G"���?D           �~@������������������������       ��?W�N�@�            r@                          �?@��U���@<           ؚ@                           �?s��C@�           �@                           �?����@           @{@������������������������       �wq��ű@�            @l@������������������������       ���?�@�            @j@                           @�j����@�           D�@������������������������       �_/�-J	@�           ��@������������������������       �s<���@           �y@                            �?I��%ȥ
@B            @\@                           @C��@             =@������������������������       ��Hַ� @
             1@������������������������       �\<����@             (@                           �?wP �%�	@0             U@������������������������       ��H8s|j	@             J@������������������������       �n{�,��@             @@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @s@     H�@      4@      K@     �{@     @T@     �@     @l@     `�@     �v@     �@@      (@     �]@     �s@      @      3@      i@      @@     h�@     �X@     �~@      e@      2@      (@     �M@     @]@      @      &@      ]@      (@     �`@     �N@      e@      W@      $@      �?      &@      A@                      :@      �?      E@      &@     �J@      3@                      @      *@                      &@      �?      9@       @      =@      @              �?      @      5@                      .@              1@      "@      8@      (@              &@      H@     �T@      @      &@     �V@      &@     @W@      I@     �\@     @R@      $@      "@      B@     �H@      @      @     @R@      "@     @R@      E@     �T@      O@      $@       @      (@      A@      �?      @      1@       @      4@       @     �@@      &@                     �M@     �h@       @       @     @U@      4@     0�@     �B@      t@     @S@       @              B@     @[@               @     �D@      2@     `j@      ?@     @_@      B@      @              1@      L@               @      <@       @     �Z@      :@     �Q@      5@                      3@     �J@                      *@      $@      Z@      @     �K@      .@      @              7@     �V@       @      @      F@       @     0w@      @     `h@     �D@      @              (@     �E@      �?      �?      :@             @p@      �?     �_@      9@                      &@     �G@      �?      @      2@       @     �[@      @     @Q@      0@      @      "@     �g@     �m@      *@     �A@     �m@     �H@     �s@      `@     @r@     �h@      .@      @     �e@      l@      &@      <@      l@     �D@     `s@     @\@     pq@     �f@      (@              H@      Q@      �?      �?     �F@      @      \@      3@     @Y@     �@@      @              8@      >@      �?      �?      6@      �?      P@      (@      H@      7@                      8@      C@                      7@      @      H@      @     �J@      $@      @      @     @_@     �c@      $@      ;@     �f@      B@     �h@     �W@     @f@     �b@      "@      @      X@     @\@      @      3@      _@      >@     @U@     @T@     �W@      X@       @              =@      F@      @       @      L@      @     @\@      *@     �T@     �J@      �?      @      1@      (@       @      @      ,@       @      @      .@      *@      .@      @              @      @                      �?      �?       @      $@      �?       @      @               @      @                              �?      �?       @              �?                       @      �?                      �?              �?       @      �?      �?      @      @      *@      @       @      @      *@      @       @      @      (@      *@              @       @      @       @      @      @      @              @      @       @                      @                              $@      @       @       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Q�ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�l�xtM@�	           ��@       	                    �?�(����@R           �@                          �<@�\mݩ@�           ��@                           �?Y�cjZ@\           Ѐ@������������������������       �(�^n^�@�            �p@������������������������       �Gn�R�@�             q@                          �>@n�S��D@'            �M@������������������������       �.�ޡ�S@             ;@������������������������       �(-QX�=@             @@
                          �9@=����B	@�           ��@                          �3@h@��v�@�           ��@������������������������       �FQ���@$           P~@������������������������       �>{W�@�           8�@                           @v�Ē��	@�            pw@������������������������       �(�&k�H	@�            �m@������������������������       �@�:��@Z             a@                           @{'���%@M           D�@                           @�����@           @�@                            �?|�F��~@           �y@������������������������       ����P9x@K             ]@������������������������       �'�"!W@�            �r@                          �4@���Q @�           ��@������������������������       �HE�V� @+           P~@������������������������       ���TUj�@�            �t@                           �?XFxܝH@E           �@                           �?����ؖ@~            �g@������������������������       ���V�s@J            �\@������������������������       �u�d�0@4             S@                          �5@���8<@�             t@������������������������       �VN�A�u@m            �f@������������������������       ��z�5��@Z            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �t@     Ȁ@      <@     �O@     �~@     �S@     P�@     �j@     8�@     �v@      4@      0@     �m@     �r@      3@     �G@     �t@     �L@     `v@     `f@     �v@     �n@      1@      �?      M@     @S@       @       @     �R@      @     `a@     �@@     `a@     �M@       @      �?      J@     �Q@       @      @     �M@      @     @a@      :@     �`@     �F@      �?      �?      7@      =@       @      @      @@      @     �S@      0@     �K@      4@                      =@      E@                      ;@              N@      $@     �S@      9@      �?              @      @              @      .@              �?      @      @      ,@      �?               @      @              @      @              �?              @      "@      �?              @      �?                      (@                      @      @      @              .@     �f@     �k@      1@     �C@     p@      J@     `k@     @b@     �k@     `g@      .@      @     `a@     �e@      ,@      A@      l@      8@     �g@      Y@      e@     @\@       @      @      E@      K@              &@     �P@      "@      ]@     �F@      T@      K@      @      @     @X@     �]@      ,@      7@     �c@      .@     �R@     �K@     @V@     �M@      @       @      E@     �H@      @      @      @@      <@      <@      G@     �J@     �R@      @      @      >@     �D@       @      @      3@      6@      (@     �A@      9@     �D@      @      @      (@       @      �?       @      *@      @      0@      &@      <@     �@@      @             @V@     �m@      "@      0@     �c@      6@      �@     �A@     �y@      ]@      @              K@      f@      �?      @     �Y@      &@     �~@      6@     �r@     �Q@       @              :@     @R@              �?     �@@       @     �a@      "@     �U@     �A@      �?               @      4@                      @             �E@      @      4@      .@                      2@     �J@              �?      >@       @     @X@       @     �P@      4@      �?              <@      Z@      �?      @     �Q@      @     �u@      *@     @j@      B@      �?              *@     �E@      �?      @      <@             �o@      @     �\@      5@                      .@     �N@                      E@      @      X@      @     �W@      .@      �?             �A@      O@       @      (@     �K@      &@      c@      *@     �]@     �F@      �?              @      <@      �?      @      (@             �P@      @      J@      0@                      @      2@              @      @             �G@              :@      "@                              $@      �?              @              4@      @      :@      @                      >@      A@      @       @     �E@      &@     �U@      @     �P@      =@      �?              &@      ,@      @      @      :@      @     �P@       @      C@      "@      �?              3@      4@      �?       @      1@       @      4@      @      <@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJq�2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��n�\@�	           ��@       	                    �?V��&T	@{           
�@                           �?�X6S��@�           ȃ@                          �;@g���f�@�            �r@������������������������       ����L@�             q@������������������������       �������@             <@                          �5@��L�@�            �t@������������������������       ��o�]�@y            �g@������������������������       ��<�>@b            �a@
                            �?��1�A�	@�           0�@                           @�#N	@            �{@������������������������       �������@           �z@������������������������       ��r�u�@
             ,@                           �?�qZ^~�	@�           L�@������������������������       ���h��	@           ��@������������������������       ���V�M@�            �q@                           @:�38��@1           �@                           �?3�O{f�@�           ��@                            �?������?�            �y@������������������������       �z헫�G�?:            �X@������������������������       �.��\
��?�            Ps@                           @����@�           (�@������������������������       ���;�@�            `n@������������������������       �?�r��@[           ��@                            �?f&���@G           8�@                           �?k��M#�@H            @^@������������������������       �ZX�j|@%            @P@������������������������       ��\���8@#             L@                           �?��dA5F@�            �x@������������������������       ��;?w�@}            �h@������������������������       �9�=
�)@�            @i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @r@     Ѐ@      <@      P@     �{@     �S@     �@     �j@     Ј@     x@      @@      4@      k@     �r@      5@     �I@     pr@      O@     �v@     �e@     �w@     �p@      <@      �?     �O@     �S@      �?      *@     �R@      @     �c@      @@      b@      L@      @      �?      =@      E@      �?       @      C@      @     @W@      0@      D@      9@      �?              9@      C@      �?      @      >@      @      W@      ,@     �C@      5@      �?      �?      @      @              @       @              �?       @      �?      @                      A@      B@              @     �B@      �?     �P@      0@      Z@      ?@      @              0@      4@              @      ,@              H@      @     �P@      3@                      2@      0@              �?      7@      �?      2@      *@     �B@      (@      @      3@      c@     @k@      4@      C@     �k@     �K@      j@     �a@     �m@     `j@      8@      �?     �D@      J@              (@     �P@      1@     �O@     �J@     �P@     �M@      $@      �?     �C@     �I@              (@     �P@      1@      O@     �G@     �P@      M@      @               @      �?                                      �?      @              �?      @      2@      \@     �d@      4@      :@      c@      C@      b@     �V@     �e@      c@      ,@      2@      V@     �]@      2@      2@      ]@      7@     �X@     �P@     �]@      _@      ,@              8@      H@       @       @     �B@      .@      G@      8@      K@      <@              �?      S@     @n@      @      *@     �b@      1@     p�@      D@     �y@     �]@      @      �?      H@      e@      @      @     �W@      @     �@      4@     r@      Q@      @              .@      H@                      3@       @     �k@       @      V@      *@                               @                      @              P@              .@      "@                      .@      D@                      0@       @     �c@       @     @R@      @              �?     �@@      ^@      @      @     �R@      @     �q@      2@      i@     �K@      @      �?      0@     �E@      �?              ;@      @     �R@      &@      F@      2@      @              1@     @S@      @      @      H@             `j@      @     �c@     �B@                      <@     �R@       @      "@     �K@      $@     �b@      4@     �^@      I@      �?              @      "@                      $@      @     �F@      @      @@      &@                       @      "@                      @      �?      5@       @      3@      @                      �?                              @      @      8@      @      *@      @                      9@     @P@       @      "@     �F@      @     �Y@      ,@     �V@     �C@      �?              "@      B@      �?      @      >@      @      J@      @     �D@      *@                      0@      =@      �?       @      .@       @     �I@      $@     �H@      :@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ#�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @+ܗ��t@�	           ��@       	                   �;@��&�>�@�           `�@                          �5@�UTev@�           ��@                           �?������@�           �@������������������������       �	�p~�@           �z@������������������������       ����IxW@�           ��@                           �?صN��@           ؈@������������������������       ����5O�@�            �q@������������������������       �><���@S           �@
                          �@@J���:q	@�             u@                           @*�y%,	@�            s@������������������������       ��[��	@�            �j@������������������������       ����k�;@3            �V@������������������������       �(W�@             ?@                           �?:�[8�g@'           d�@                          �4@i~�$@@`           ��@                           �?�ph��?�            �u@������������������������       �^���i�?t             h@������������������������       �^.�Rҧ�?`            �b@                           @?����@�            `k@������������������������       �{~���@B             Y@������������������������       ��&w�z�@J            �]@                          �4@ ��k�@�           ��@                           @F�k @b            �@������������������������       ��5���D@R            �`@������������������������       ����-@           �y@                           @Z-t�G @e           0�@������������������������       ���p�t�@X           ��@������������������������       �}r%RFS@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@     �s@     0�@      B@      M@     �|@     �S@      �@     �j@     @�@     �u@     �@@      3@     @l@     0u@      7@     �F@     Pt@     �M@     x@      f@      w@      m@      ;@      "@     �g@     �q@      4@     �@@     �q@     �G@     �v@      a@     �t@     �d@      9@      "@     @X@     �b@      "@      0@     @c@      4@     �o@     �Q@     �j@      V@      $@      @     �C@     �N@      "@      @     @R@      "@     �Z@      ?@     �O@      :@       @      @      M@     �V@              $@     @T@      &@     `b@     �C@      c@      O@       @             �V@     �`@      &@      1@     �`@      ;@      [@     �P@      ]@     @S@      .@              A@     �H@      �?      *@      F@      @     �F@      0@     �L@      0@      @             �L@     �U@      $@      @      V@      8@     �O@      I@     �M@     �N@      "@      $@      C@     �J@      @      (@     �C@      (@      7@      D@     �B@     �P@       @      @     �@@      J@      @      (@      >@      &@      6@      A@     �B@      P@       @      @      7@      H@      @      "@      4@      @      &@      9@      ;@     �B@       @              $@      @              @      $@      @      &@      "@      $@      ;@              @      @      �?                      "@      �?      �?      @              @              �?     @V@     `n@      *@      *@      a@      4@     ��@      C@     �y@     �\@      @              .@     @U@       @      �?      6@      @     �p@       @     �`@      7@       @               @      D@              �?      (@             �g@      @      R@      *@       @              @      3@              �?      &@              ]@      @      <@      $@                      @      5@                      �?             �R@       @      F@      @       @              @     �F@       @              $@      @     �R@      @     �N@      $@                      @      4@                      @      @     �D@              2@      @                      @      9@       @              @              A@      @     �E@      @              �?     �R@     �c@      &@      (@     �\@      ,@     Pu@      >@     0q@      W@      @              =@     �S@      @       @      B@       @     @k@      &@     �`@      ?@                      .@      =@                      "@       @      F@      @      7@      @                      ,@     �H@      @       @      ;@             �e@      @     @[@      9@              �?     �F@      T@      @      $@     �S@      (@     �^@      3@     �a@     �N@      @      �?     �B@     �S@      @      $@     �R@      "@     �^@      3@     �a@     �N@      @               @      �?      @              @      @      �?              �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ahG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              �?e��qU@�	           ��@                           @)���y�@�           ��@                           @*�֗$@�           ؅@                           �?�d�@�           X�@������������������������       ����BL�@�            0p@������������������������       �'֎}�@            �z@������������������������       �|R��>@	             0@                           �?��L@�             x@	       
                    �??��ԏL @N            �_@������������������������       �QN�� ��?%             P@������������������������       ��@hi� @)             O@                           �?�Ǣ@�            @p@������������������������       ����0<�@V            @`@������������������������       ���\��b@Q            @`@                           �?���mh@           �@                           �?u�bns@9           ��@                          �8@��7�P@�            �t@������������������������       � mgj�@�            �o@������������������������       �d�(e�@3            �S@                            @T_��@a           X�@������������������������       �_�(=Y@           �y@������������������������       ���)�L�?Y            �a@                           @�+ae]T@�           X�@                           @A��	@�           �@������������������������       �<�T�	�	@j           h�@������������������������       ���aA8	@O            �^@                            @t��y�@+           x�@������������������������       ���A�1@�           ��@������������������������       ��x�lRJ@v            @g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     @s@     0�@      A@      L@      z@     �T@     ��@      i@     ��@     �u@     �D@       @      T@     �b@              5@     �\@      2@     �r@     �K@     �k@      [@      2@       @      O@     �W@              3@     �W@      *@     @a@     �D@     `a@     �S@      2@       @      M@      W@              3@      W@      *@     @a@      D@     `a@     �S@      (@       @      7@     �F@              @      G@      @      I@      3@      G@      .@      @             �A@     �G@              0@      G@       @      V@      5@     @W@     �O@      @              @       @                       @                      �?              �?      @              2@      L@               @      4@      @     �c@      ,@      U@      =@                              7@                      @      @     �O@       @      7@      @                              $@                      @      �?     �@@              *@      @                              *@                      @       @      >@       @      $@       @                      2@     �@@               @      ,@       @     �W@      (@     �N@      7@                      @      4@               @      *@             �C@      @      ?@      (@                      &@      *@                      �?       @      L@      @      >@      &@              0@     �l@      {@      A@     �A@      s@     @P@     P�@     @b@     ��@     �m@      7@             �S@     �]@      @      @     �R@      @     t@      ;@     �h@      H@      @              F@      M@      @      @     �F@       @     �Q@      1@      J@      ?@      @             �@@      G@      @              8@       @     �O@      0@     �E@      5@      �?              &@      (@              @      5@               @      �?      "@      $@       @             �A@     �N@               @      =@      @     @o@      $@     `b@      1@      �?              >@      J@                      5@      @      f@      "@     �Z@      .@      �?              @      "@               @       @             @R@      �?     �D@       @              0@     �b@     �s@      >@      =@     �l@      N@     �x@     �]@     �x@     �g@      3@      .@     �Y@      g@      9@      2@     @c@     �H@     �`@     �X@     �d@     �`@      0@      $@     @W@     �d@      9@      2@     �`@      E@     @\@     @U@     �c@      _@      "@      @      "@      4@                      6@      @      4@      ,@       @      $@      @      �?     �G@      `@      @      &@      S@      &@     @p@      4@     �l@      K@      @      �?      F@     �Z@      @      "@      J@      $@      h@      ,@     �f@      G@      @              @      5@       @       @      8@      �?      Q@      @     �I@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ")ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @�kn��@�	           ��@       	                     �?�m$.�@j           ڠ@                           �?�����)@�           ؅@                          �;@?���@�            @j@������������������������       ���n=u
@x            �g@������������������������       ��v+��s@             6@                          �2@$�AF!�@0           �~@������������������������       ��4a���@8             X@������������������������       ���)�	@�            �x@
                          �2@�����@�           Ȗ@                           �?g�ǎ�@�            @t@������������������������       ��-���@�            �n@������������������������       �M�|��@9             T@                           �?��E�nI	@�           ��@������������������������       ��d����@�            �r@������������������������       �M�}�	@           (�@                          �4@��ǶC�@Q           p�@                           @�ݣ��@R           �@                          �1@J* C�� @�           ��@������������������������       ��lw��V�?�             q@������������������������       ���H�@�            pv@                           �?_���@�            �t@������������������������       ���u`Ѫ@^            @c@������������������������       �PR���r @i             f@                           @����@�           Ј@                           @f��K)�@�           0�@������������������������       ���<�~8@F           �@������������������������       ��.Xm�d@�            �p@������������������������       ���L��( @	             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     �q@     ��@      =@     �G@     p}@     �U@     ��@     @k@     h�@     `t@     �@@      2@     @h@     �s@      3@     �@@     �t@     @P@     �w@     `f@     �x@     �i@      <@      @     �M@     �W@       @      &@     �X@      6@      a@      P@     �b@     �E@      ,@      @      3@      @@               @      .@      �?     �J@      @     @Q@      $@      �?              1@      >@               @      (@             �J@      @      P@      @              @       @       @                      @      �?                      @      @      �?              D@      O@       @      "@     �T@      5@      U@      N@     �T@     �@@      *@              @      4@                      *@      @      >@      @      1@      @                     �B@      E@       @      "@     �Q@      2@      K@      K@     @P@      =@      *@      ,@     �`@     @k@      1@      6@      m@     �E@     �m@     �\@     �n@     @d@      ,@      �?      1@      F@                      K@       @     �U@      3@      O@      B@       @      �?      &@      B@                     �G@       @     �L@      (@      G@      >@       @              @       @                      @              >@      @      0@      @              *@     �]@     �e@      1@      6@     `f@     �D@      c@      X@      g@     �_@      (@              A@     �A@      �?      @     �E@             �P@      5@     �N@      <@       @      *@      U@     `a@      0@      1@      a@     �D@     @U@     �R@     �^@     �X@      $@      �?     @V@     �k@      $@      ,@     �a@      5@     @�@     �C@      z@     @^@      @             �@@     �\@      @      $@     �J@      @     �{@      $@      n@      I@      �?              8@     �S@      @      @     �A@       @     �s@      @     �a@      2@      �?              (@      9@              �?      1@              d@             �I@      @      �?              (@     �J@      @      @      2@       @     �c@      @     �V@      *@                      "@     �B@              @      2@      @      _@      @     �X@      @@                       @      .@              @      ,@             �N@      @     �A@      (@                      �?      6@                      @      @     �O@              P@      4@              �?      L@     @Z@      @      @     �U@      0@     �m@      =@     �e@     �Q@      @      �?     �G@     @Z@      @      @     �U@      $@     �m@      ;@     �e@     �Q@      @      �?      =@     �Q@              �?     �H@      @     �f@      .@     �\@     �A@      @              2@     �A@      @      @     �B@      @     �K@      (@      N@      B@      �?              "@              �?              �?      @      �?       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJy��`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @_e���!@�	           ��@       	                    �?�����@Y           �@                           �? ���	@�           �@                           �?����@            �@������������������������       �����?@�            p@������������������������       ����-�@�            0v@                           �?"��7ϛ	@v           �@������������������������       �9 �TV@�            Pq@������������������������       ����3Q"
@�           @�@
                            @V��@�@d           ��@                          �=@`����@           �y@������������������������       ���.�[k@�            0x@������������������������       ��˨�ڒ@             9@                           �?����@^            �c@������������������������       ���O>��@*             R@������������������������       ��g�1�|@4             U@                          �4@ZS�*�@W           @�@                           �?-����@]           �@                           �?:-�@>           �~@������������������������       ��_B��K�?�             l@������������������������       �L�u���@�            �p@                           @=�+i@           p{@������������������������       ���� ��@Q            �_@������������������������       ��oG?�@�            �s@                           @�}�k^�@�           p�@                           @��3;Z@�           Ȉ@������������������������       �Y� �@:           `@������������������������       ���z��@�            0r@                          �8@��#Qw#@             5@������������������������       �QcX^@             $@������������������������       �=*,I�R @             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     H�@      ?@      P@     �y@     @U@     А@     �h@     ��@     v@      ;@      ,@     �l@      u@      3@     �G@     �p@     �M@      x@      d@     �w@      o@      7@      ,@     @g@      n@      1@     �D@      i@      D@     `n@     �^@     �p@     `i@      6@      @     �J@     �V@      �?      (@      T@      $@      _@      @@     �^@     �R@      "@      @      0@     �J@              @      C@      @     �K@      "@     �E@      <@      @             �B@      C@      �?       @      E@      @     @Q@      7@     �S@     �G@      @      &@     �`@     �b@      0@      =@     @^@      >@     �]@     �V@     �b@      `@      *@              D@     �H@      �?      @      :@      @      G@      3@     �J@     �@@              &@     @W@     @Y@      .@      6@     �W@      ;@     @R@     �Q@      X@     �W@      *@              F@     �W@       @      @     @P@      3@     �a@     �C@     �[@     �F@      �?             �A@     �L@       @      @      I@      .@     �W@      @@     �W@      <@      �?              8@     �L@       @       @      G@      *@     @W@      <@     �W@      <@                      &@                      �?      @       @       @      @                      �?              "@      C@              @      .@      @      G@      @      1@      1@                      @      &@                      @      @      7@      @      (@       @                      @      ;@              @      "@              7@      @      @      "@              �?     �T@      k@      (@      1@     �a@      :@     ��@     �A@     �y@     @Z@      @              @@     �Z@      @      &@      M@       @     �{@      (@     @j@      H@      �?              (@     �I@      @       @     �A@      @      o@       @     �X@      8@                      @      6@              @      @             �a@      �?     �B@       @                      @      =@      @      @      >@      @     @Z@      @      O@      0@                      4@     �K@              @      7@      @      h@      @     �[@      8@      �?               @      :@                       @      @     �K@              8@      @                      (@      =@              @      5@             @a@      @     �U@      2@      �?      �?     �I@     �[@      "@      @     @U@      2@     `o@      7@     �h@     �L@      @      �?     �G@     @[@       @      @     @S@      ,@     `o@      6@     �h@     �L@      @      �?     �A@      Q@              @     �E@       @     @g@      @     �]@      =@      @              (@     �D@       @      @      A@      @     @P@      .@     �S@      <@                      @       @      �?               @      @              �?      �?                               @              �?              @      @              �?                                       @       @                      @      �?                      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJM��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\��      C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��ČD@�	           ��@       	                   �8@�u�l�@�           ��@                           �?����4@�           �@                            @�i��@8           �~@������������������������       �Ulڜr�@�            �r@������������������������       �����I@s            �g@                          �4@G�����@�           L�@������������������������       �����y{@y           ��@������������������������       �ef���@@           p@
                            @pu����	@�           0�@                            �?��kY�@�            �x@������������������������       ��F�8"1	@�            �s@������������������������       �820d!@,            @U@                          �=@0`���O
@�             o@������������������������       �JѰ8I
@k            �d@������������������������       ��O��D)@,            �T@                          �6@�e��.�@"            �@                           @��C�	@�           @�@                           �?w:��F�@�            p@������������������������       ���ڞ@P             _@������������������������       �\�5��^@S            �`@                           �?�o�H@=           x�@������������������������       �8�-����?�            �t@������������������������       � �(�)@l           (�@                          �8@�����A@B           �@                           @�i���@�             k@������������������������       �}<?I�@            �D@������������������������       �7樖n�@m            �e@                           �?"u��\�@�             r@������������������������       ��d�5�P@O             `@������������������������       �KMٲ(#@l            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �s@     ��@     �@@      J@     �{@      T@     ؎@      i@     ȉ@     �v@      :@      1@      m@     �u@      :@      F@     �r@      P@     �v@     �c@     �x@     �p@      :@       @     �c@     @o@      .@      @@     �i@      C@      r@      Y@     �t@     `c@      *@             �K@     �R@      �?      @     �D@       @     @`@      7@     �]@     �B@       @              C@      B@      �?      @      :@      �?     @T@      ,@     @S@      3@       @              1@      C@              �?      .@      �?     �H@      "@      E@      2@               @     �Y@      f@      ,@      <@     �d@      B@      d@     @S@     @j@     �]@      &@      @      B@     �U@      "@      "@      V@      *@     @Z@      J@     �^@     �Q@       @      @     �P@     �V@      @      3@     �S@      7@     �K@      9@      V@     �G@      @      "@     �R@     �X@      &@      (@      X@      :@      R@     �M@     �P@     @[@      *@      @      E@     �J@      @       @     �P@      ,@      F@     �A@      F@     �S@       @       @      A@     �F@      @       @      E@      *@      B@     �A@     �@@      M@       @      @       @       @                      9@      �?       @              &@      4@              @     �@@     �F@      @      $@      =@      (@      <@      8@      6@      ?@      @      �?      7@      3@      @      @      5@      (@      2@      5@      4@      3@      @       @      $@      :@      @      @       @              $@      @       @      (@              @      T@     �k@      @       @     @a@      0@     ��@      E@     �z@     �Y@                     �B@     �d@      @      @     �S@       @     0@      0@     �r@      N@                      2@      G@                      0@      @     @X@      @     �J@      *@                      (@      *@                      &@      @     �F@      @      6@      &@                      @     �@@                      @       @      J@       @      ?@       @                      3@      ^@      @      @      O@      �?      y@      "@     `n@     �G@                      @      E@              �?      1@             �g@      @     @P@      @                      (@     �S@      @       @     �F@      �?     �j@      @     @f@      E@              @     �E@      K@       @      @      N@       @     �_@      :@     �`@     �E@              @      <@      =@      �?      �?      ;@      @     �J@      @      K@      *@              @              @                      �?      �?      *@              .@      @                      <@      9@      �?      �?      :@       @      D@      @     �C@      "@                      .@      9@      �?      @     �@@      @     @R@      6@      T@      >@                      @      1@              �?      *@              F@      (@      =@      @                      "@       @      �?      @      4@      @      =@      $@     �I@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJPq�
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�b��@@�	           ��@       	                   �7@� ��!�@r           4�@                          �5@��}*�@�           ��@                           �?g4�u@�           ��@������������������������       ��9� ��@�            �x@������������������������       �C�	Zz@�           ��@                           @�̚�@�            @t@������������������������       ��;i�@t             f@������������������������       ��E�1#?@_            `b@
                          �<@��f��	@�           ��@                           �?��Ȭ	@I           �@������������������������       ��J~�6@[            �`@������������������������       ���F�	@�            0w@                          @@@���z}F	@�            `o@������������������������       �*Āv�4	@|            �i@������������������������       �����k@            �G@                           @0ATFl"@G           ��@                          �4@yj�U*@�           x�@                           �?6���=@�           p�@������������������������       �_^ a�@�            �u@������������������������       ��%�`}e @�            0u@                           @�;e�~�@H            @������������������������       �-u�'eq@>           0~@������������������������       �GC7�K@
             *@                           �?�%7�@K           ��@                          �0@C�����@~             i@������������������������       ��K�Qp� @             3@������������������������       ��C�6-@s            �f@                          �5@�-0�~n@�            �t@������������������������       ��c	�l/@k            @e@������������������������       �K����@b            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     �@     �@@     �J@     �|@     �S@     ��@     @j@     ��@     �u@      ?@      0@     �k@     �s@      =@     �A@     pt@     �M@     @y@     `d@     �v@     `n@      :@      $@     �b@     �i@      "@      7@      j@      5@     �s@     �U@     �p@      a@      (@       @     �W@     @b@       @      *@     �c@      3@     �p@     �Q@     �l@      Z@      @              @@     �H@                     �B@      @      _@      1@     �Y@      >@      �?       @     �O@     @X@       @      *@     �^@      0@     �a@     �J@     @_@     �R@      @       @     �K@      N@      �?      $@     �H@       @      H@      0@     �E@     �@@      @      �?      ;@      :@      �?      @      <@             �B@      @      <@      4@              �?      <@      A@              @      5@       @      &@      (@      .@      *@      @      @     �Q@     �[@      4@      (@     �]@      C@     �V@     @S@      W@     �Z@      ,@      @     �J@     �R@      .@      @     �R@      1@     �R@     �H@     �Q@     �L@      (@      �?       @      2@                      7@              <@      *@      .@      6@      @       @     �F@      L@      .@      @     �I@      1@      G@      B@     �K@     �A@      @      @      2@      B@      @      @     �F@      5@      1@      <@      6@     �H@       @       @      ,@      ?@       @      @     �@@      4@      1@      9@      ,@     �C@       @      �?      @      @      @              (@      �?              @       @      $@              �?     �S@     Pp@      @      2@     �`@      4@     ��@     �G@     @{@     �Y@      @      �?      K@     �g@              @     @T@      $@     �{@      9@     @s@      N@      @              9@     �[@               @      :@       @     `r@      (@     @g@      =@                      1@      M@                      1@             �a@       @     @V@      1@                       @      J@               @      "@       @      c@      @     @X@      (@              �?      =@     @T@              �?     �K@       @      c@      *@     �^@      ?@      @      �?      ;@     @T@              �?     �I@      @     �b@      "@     �^@      ?@      @               @                              @       @      �?      @                                      8@     �Q@      @      .@      J@      $@      d@      6@      `@      E@       @              @      >@      �?      �?      3@             �R@      @     �K@      (@                               @                      @              @              �?      @                      @      6@      �?      �?      .@             �Q@      @      K@      "@                      5@      D@      @      ,@     �@@      $@     �U@      0@     @R@      >@       @              @      :@              @      *@       @     @P@       @     �B@      (@       @              .@      ,@      @      "@      4@       @      5@      ,@      B@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ)6F4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@6����5@�	           ��@       	                    �?T��Hp�@�           ��@                           �?]�����@�            �v@                           �?�����@\            `c@������������������������       ��f���b@.            @T@������������������������       ��8^�A�@.            �R@                          �0@��\�D@�            `j@������������������������       ��+��[@             @@������������������������       ��
!,�@r            `f@
                           @�C�J(@�           ��@                          �1@f6���V @c           ؁@������������������������       �ֽ�$G-�?�            �u@������������������������       �횊�r@�             l@                          �0@�_�v�@\            ``@������������������������       ���״�1@             3@������������������������       ��ҏ��d@N             \@                          �<@����@           :�@                           �?n��A�@?           ��@                          �9@1Itd!@�           @�@������������������������       �
M߂@�           ��@������������������������       �j^�z��@E            �\@                          �5@޿g��g@o           X�@������������������������       ��-�E�@�           ��@������������������������       �� �@q           0�@                            �?�0`S5	@�            �s@                          �=@��}�A@j            �d@������������������������       �^�b^x�@&            �N@������������������������       ��8��@D            @Z@                           �?�r����@^             c@������������������������       �<sx8V@            �E@������������������������       ����<@B            �[@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     s@     �@      :@     �P@     �}@     �R@      �@     �h@     ��@     u@      <@      @      M@     �_@       @      @      \@      �?     @z@      ?@     �m@      P@      @      @      @@     �H@              @     @Q@      �?     �T@      6@     @Q@      ?@      @      @      &@      3@                      A@      �?     �E@      "@      .@      0@       @       @      @      &@                      2@      �?      =@      �?      @       @              @      @       @                      0@              ,@       @      $@       @       @              5@      >@              @     �A@             �C@      *@      K@      .@      �?              @      "@              �?       @              "@       @      �?       @                      .@      5@               @     �@@              >@      &@     �J@      *@      �?              :@     @S@       @      @     �E@              u@      "@      e@     �@@       @              4@     �P@       @      �?      =@             0r@      @     ``@      7@                      $@      >@                      *@             @h@      @     @U@      (@                      $@     �B@       @      �?      0@             @X@      @      G@      &@                      @      $@               @      ,@             �G@       @      C@      $@       @                      @                      �?              @              @      @                      @      @               @      *@             �D@       @     �@@      @       @      2@     �n@     �y@      8@      N@     �v@     �R@     ��@     �d@      �@     q@      7@      0@      j@     �w@      5@      I@     Ps@     �L@     ��@     �a@     (�@     �i@      3@              L@     @]@      @       @     �P@      "@     �i@      1@      g@      D@       @             �I@      V@      @       @     �I@      @     �f@      .@     `c@     �C@       @              @      =@                      0@      @      9@       @      >@      �?              0@      c@     0p@      1@      E@     @n@      H@     �v@     �^@     �v@     �d@      1@      @     �E@     �\@      @      .@     �\@      4@     @h@     �H@     `e@      S@      @      $@     @[@      b@      $@      ;@     �_@      <@     �e@     �R@      h@     �V@      (@       @     �C@     �C@      @      $@      J@      1@      >@      :@      ?@     �P@      @      �?      1@      3@              �?      3@      (@      (@      3@      2@      F@      @      �?      @      $@              �?      @      @      @      @      @      ;@                      ,@      "@                      ,@      "@      "@      0@      *@      1@      @      �?      6@      4@      @      "@     �@@      @      2@      @      *@      6@                              "@              @      @              *@      �?      @      @              �?      6@      &@      @      @      ;@      @      @      @      @      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�@�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��$�@�	           ��@       	                   �:@"�.�z�@�           ��@                          �4@�$
�@@�           ��@                           �?P� .v�@2           �@������������������������       ��;�@�           ȃ@������������������������       ��LH=�@�            �p@                           �?���{hD@N           (�@������������������������       �)vJ��@�            �q@������������������������       ���tQ�@�           @�@
                           �?U����
@            {@                          @@@,����	@�            Pv@������������������������       ��>��N�	@�             s@������������������������       �٩���@!            �I@                          �<@�H��u2@2            �R@������������������������       ���U��@            �A@������������������������       ��'(��@             D@                           @��:+�i@(           ̙@                            @����@�           ��@                           @��1CL�@8           ��@������������������������       �{!w:�@Q           ��@������������������������       �}呴@�            @u@                           @<�*C�=@�            @o@������������������������       �&z�7G@H            �\@������������������������       �Y��@N             a@                           @��i���@Z            `b@                            �?��s�թ@F             [@������������������������       ���d@V@%            �N@������������������������       �-�u憹@!            �G@                           7@ɰ���H	@            �C@������������������������       �V@���@             *@������������������������       �IW����@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �t@     ��@      >@      N@     @@     �T@     ��@     �l@     ��@     �u@      C@      1@      n@      u@      4@     �F@     Pv@     �N@     w@     �g@     @v@     @n@      <@      @      h@     Pr@      .@     �A@     �q@     �D@     �t@     @a@     �s@     @d@      1@      @      M@      _@      &@      (@     �a@      &@      h@     �R@     �d@     �W@       @      @     �D@     @T@      @      "@     �[@      &@      \@     �J@      ^@     �S@       @              1@     �E@      @      @      @@              T@      6@     �F@      0@              �?     �`@      e@      @      7@      b@      >@     �a@     �O@     �b@     �P@      "@              H@      G@      �?      @      ;@      @     �P@      &@      Q@      $@       @      �?     �U@     �^@      @      4@     �]@      ;@     �R@      J@      T@     �L@      @      (@      H@     �F@      @      $@     �Q@      4@     �B@     �I@     �E@      T@      &@      (@      E@      A@      @      "@     �M@      0@      6@      D@      A@     �R@      $@      &@     �A@      <@       @      @     �I@      0@      5@     �B@      6@     �P@      $@      �?      @      @      @       @       @              �?      @      (@       @                      @      &@              �?      &@      @      .@      &@      "@      @      �?              @      @                      @              (@      @      @      �?                      @      @              �?      @      @      @       @      @      @      �?             �W@     �i@      $@      .@     �a@      5@     �@     �C@     �x@     @Z@      $@             @R@     @h@      @      ,@     @`@      3@      �@      =@     @w@      W@       @             @P@      g@      @      "@      [@      ,@     0}@      :@      s@      R@       @             �E@     @a@              �?     �Q@      "@      x@      .@      i@     �J@      �?              6@      G@      @       @      C@      @     �T@      &@      Z@      3@      �?               @      $@              @      6@      @     @[@      @      Q@      4@                      @      @              @      @      @     �O@      @      6@      @                      @      @               @      0@       @      G@              G@      0@                      5@      &@      @      �?      *@       @     �A@      $@      :@      *@       @              (@       @       @              $@      �?     �@@      @      5@      (@      @              "@      @       @                      �?      9@       @      &@      @                      @      @                      $@               @      @      $@      @      @              "@      @      @      �?      @      �?       @      @      @      �?      @               @                      �?      @                              @              @              @      @      @                      �?       @      @       @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ� "thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�Ah=�B@�	           ��@       	                   �8@D;C�@e           ֠@                          �1@�s�F�Q@�           H�@                          �0@�!��j�@�            `q@������������������������       ��8�@:             V@������������������������       �[&���@v            �g@                            @�~�W�@3           �@������������������������       �3Z��@�           ��@������������������������       ���b\L@5           @~@
                           �?W#�s�v	@�           Ȃ@                           �?�3���@�            �n@������������������������       �������@8             X@������������������������       ���ň�@a            �b@                          �:@��Y�&�	@�            @v@������������������������       ��ePKc@Q            �^@������������������������       �L�
y	@�            @m@                           @1�@K           x�@                          �2@S��w�@�           �@                            �?��u*X�?           p{@������������������������       ���?ս�?>             Y@������������������������       �KIR� @�            0u@                           @�J!(@�           h�@������������������������       �>٬��@;           �@������������������������       �伞4Rh@�            Pq@                          �5@w�8@U           Ѐ@                          �3@���$�.@�            @s@������������������������       �G�|�n@�            �h@������������������������       ���-�@E            �[@                          �6@���d��@�            �l@������������������������       ����f�@             B@������������������������       ��9u@{            @h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@      s@      �@      B@      L@     �z@      T@     �@     �i@     ��@     �v@     �A@      *@     �k@      t@      9@     �D@     s@     �N@     �u@     �d@     �x@     �m@      <@      @     �`@     �l@      4@      >@      n@     �B@     @q@     �Y@     �s@     @b@      0@      �?      5@     �C@      �?       @     �B@              S@      0@     �N@      8@                      "@      0@               @      3@              0@      @      *@      $@              �?      (@      7@      �?              2@              N@      *@      H@      ,@              @     @\@     �g@      3@      <@     `i@     �B@      i@     �U@     �o@     �^@      0@      �?     �U@     �X@      *@      3@      ^@      7@     �_@     �N@     `d@     �Q@      $@      @      ;@      W@      @      "@     �T@      ,@     @R@      9@      W@      J@      @      @     �U@     �V@      @      &@     @P@      8@     �Q@      O@     �S@     �V@      (@      �?     �@@     �B@      @      @      >@      $@      :@      4@      @@      H@                      &@      .@               @      (@              ,@      @      1@      2@              �?      6@      6@      @      @      2@      $@      (@      *@      .@      >@              @      K@     �J@       @      @     �A@      ,@      F@      E@     �G@      E@      (@              .@      <@              @      *@      @      (@      2@      1@      @       @      @     �C@      9@       @      @      6@      $@      @@      8@      >@      C@      @      �?     �T@     �l@      &@      .@      ^@      3@     �@      E@     �z@      `@      @      �?      M@     @c@      @      @     �Q@      $@     P�@      6@     r@     �T@      @              6@      F@       @              ,@      �?      n@      @     �W@      ,@                      �?      @                       @             �R@              *@      @                      5@     �C@       @              (@      �?     �d@      @     �T@      "@              �?      B@     �[@       @      @      L@      "@     �q@      0@     @h@      Q@      @      �?      ;@      R@       @              F@      "@     @c@      ,@     @`@     �G@      @              "@      C@              @      (@             �_@       @      P@      5@                      9@     �R@      @      &@      I@      "@      c@      4@     `a@     �G@      @              &@      G@      �?       @      9@      �?     @Z@      @     �T@      4@      @              @      1@      �?      @      4@             @Q@      @     �M@      .@                      @      =@              �?      @      �?      B@       @      8@      @      @              ,@      <@      @      @      9@       @      H@      .@      L@      ;@                              �?       @               @      @      @              @      "@                      ,@      ;@      @      @      1@      @      E@      .@      I@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ弟OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?l�A�@�	           ��@       	                    @��RFp@@           ��@                           �?Ю���@�           ��@                          �;@�D(e@�            �w@������������������������       �v>�;Y@�            �t@������������������������       �6(�i8@            �F@                           @���n�a	@�           x�@������������������������       �p"��[@�             u@������������������������       ��ZT.�	@           �y@
                           �?�]��+�@n           Ȏ@                           @��`U@E           �@������������������������       �&�'W`@[            `c@������������������������       �f��c@�             v@                            �?,u�	��@)           �}@������������������������       �g&��%y@}             j@������������������������       ��N�0��@�            �p@                          �5@N��u�@f           $�@                           �?��Q�,�@c           ��@                           �?8���3@�            `v@������������������������       �5�H�@q            �g@������������������������       �HҞ_У@l            @e@                           �?����@�           ȃ@������������������������       ��f�z��@�            `o@������������������������       �e�����@�            �w@                           �?/��;O�@           P�@                           �?�rQʹf@�            �j@������������������������       ��Jb{��@L            �]@������������������������       ��_"��p@=             X@                           @��#��,@z           ��@������������������������       �?�g�G@@�            �v@������������������������       �*��&	@�            @m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        @     @s@     ��@      ;@      J@     �|@      S@     ��@     �j@     ��@      w@     �@@      @      e@     �p@      0@      A@     �l@      L@     P�@      `@     �|@     `i@      3@      @     �\@     �c@       @      :@     �a@     �G@     �f@     �W@     @j@      `@      1@       @     �E@     �H@      �?      @     �C@      �?     @T@      3@     �W@      A@      @             �A@     �E@      �?      @      A@             �S@      0@     �V@      6@      @       @       @      @              �?      @      �?       @      @      @      (@      �?      �?     �Q@     �Z@      @      4@     �Y@      G@     �Y@     �R@      ]@     �W@      $@              =@     �E@              &@     �I@      8@     �I@      3@     �M@      H@      �?      �?      E@      P@      @      "@     �I@      6@     �I@      L@     �L@      G@      "@             �K@     �\@       @       @      V@      "@     0u@      A@     �o@     �R@       @             �B@      O@              @      K@      @     �e@      &@     @`@      <@       @              6@      9@                      1@      @      J@      @      3@      &@       @              .@     �B@              @     �B@      �?     �^@      @     �[@      1@                      2@     �J@       @      �?      A@      @     �d@      7@     �^@     �G@                      "@      2@      @              "@      @     �W@      $@     �D@      .@                      "@     �A@      �?      �?      9@      �?     �Q@      *@     @T@      @@               @     `a@     �p@      &@      2@     �l@      4@     �~@      U@     @v@     �d@      ,@             �F@     �a@       @      $@     �[@      "@     `u@     �B@     �i@     �T@      @              3@     �E@               @      8@      �?     �c@       @     �T@      3@                      @      5@              �?      &@      �?     �V@      @     �D@      &@                      *@      6@              �?      *@              Q@      @      E@       @                      :@     �X@       @       @     �U@       @     �f@      =@     �^@     �O@      @              (@      C@       @      @     �B@      @     �R@      @     �D@      A@      @              ,@      N@              @      I@      @     @[@      9@     �T@      =@      @       @     �W@     @`@      "@       @     @]@      &@     �b@     �G@     �b@     @U@       @              2@      D@       @      @      1@       @     �N@      @     �I@      .@                      @      <@       @      @      $@      �?      :@       @      B@      @                      *@      (@                      @      �?     �A@      @      .@      $@               @      S@     �V@      @      @      Y@      "@      V@      E@     �X@     �Q@       @       @     �M@     @P@      @             �J@      @      @@     �@@      F@      K@       @              1@      9@       @      @     �G@      @      L@      "@     �K@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJk%qqhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�K��H@�	           ��@       	                   �<@��c�pb@/           (�@                           �?�~|O�@�           ��@                           �?Q�sܰ	@�           ��@������������������������       ��^�V�@z            `g@������������������������       �6��b�;@           @|@                          �7@�����@`           h�@������������������������       ��U�5�@           `{@������������������������       �(��i��@O            �]@
                           @�_W�}@9            �W@                          @@@Pm(;@*            �P@������������������������       �@�(��\@!            �I@������������������������       ��"�@}��?	             .@                            �?��th�@             <@������������������������       �݁N)��@             3@������������������������       �Sn�K�A�?             "@                           @�a>CBL@�           ~�@                           �?��c�%{	@�           X�@                            �?�9��y�	@�           ؐ@������������������������       �]�c��@�            �t@������������������������       �y�2N�
@�           P�@                            �?@n��pX@            z@������������������������       ��;��@G            @\@������������������������       ����Ny�@�            �r@                          �5@��hIY@�           ��@                           @�F�mF�@�           Ѕ@������������������������       ��2�(��@G           �@������������������������       ��?�"��@s             g@                          �:@����@            �z@������������������������       ������@�            `r@������������������������       �敐*��@U             a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     pr@     ��@      >@     �P@     �}@     �R@     D�@      k@     8�@     �t@      =@      �?      V@     `e@      @      &@     �^@       @     �~@     �E@     �p@     @T@      @      �?     @T@     �c@      @       @     @Z@       @     �}@      >@     @p@      M@      @      �?     �B@      V@      @       @     @Q@      @     `p@      7@     �]@      7@       @      �?      3@      6@      @      @     �@@             �D@      3@      @@      "@       @              2@     �P@               @      B@      @     �k@      @     �U@      ,@                      F@     �Q@                      B@      @      k@      @     �a@     �A@       @              C@      I@                      5@              g@      @      [@      ?@                      @      5@                      .@      @      @@       @     �@@      @       @              @      (@              @      2@              $@      *@       @      7@                      @      @              @      ,@              @      $@       @      4@                      @      @                      @              @       @      �?      4@                      �?                      @       @                       @      �?                                      @                      @              @      @      @      @                              @                      @              @      @      @      �?                              �?                                      @              @       @              4@     �i@     `x@      ;@      L@     �u@     �P@     @�@     �e@     �@     @o@      9@      3@      a@     �l@      0@     �D@     �m@      J@     �i@      c@      l@     �c@      5@      3@     �[@      c@      0@      A@     �f@      D@      ]@     @\@     `c@     �^@      3@      �?     �C@     �B@      �?      $@     �K@      "@     �B@     �H@     �M@      ;@       @      2@     �Q@      ]@      .@      8@     @_@      ?@     �S@      P@      X@      X@      &@              ;@      S@              @      L@      (@     �V@      D@     �Q@      B@       @              @      <@               @      ,@       @      <@      @      ,@      "@       @              7@      H@              @      E@      @      O@      B@      L@      ;@              �?     �Q@      d@      &@      .@     @\@      ,@     �u@      5@     �q@     �V@      @              >@     �X@      @       @      L@      @     @m@      @     �i@     �E@      @              3@      R@      �?      �?     �A@      @     `g@      @     `c@      >@      @              &@      ;@      @      @      5@       @     �G@       @      I@      *@              �?      D@      O@      @      @     �L@      @      \@      ,@     @S@      H@      �?      �?      5@      E@      @       @      ?@      @     �T@       @     �N@     �@@      �?              3@      4@      �?      @      :@              =@      @      0@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ChG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?�B��q@�	           ��@       	                    �?L�-�?�@�           ��@                           @<��R��@           @z@                          �7@o�d��O@�            Pp@������������������������       �j9eސ}@{            �g@������������������������       ������@/             R@                           @!�DG�)@e            �c@������������������������       �/s����@O            �_@������������������������       �o)	{@             @@
                          �4@F��u@y           ��@                           �?y���z@�            �p@������������������������       �q��aP�@>            �V@������������������������       ���8�� @k            �e@                           �?S�,��	@�            �t@������������������������       ��0j�Pf@1            �S@������������������������       ��i�M|	@�             p@                           @o�X$V@A           ��@                          �2@����@�           |�@                           �?�cp%�c@�             v@������������������������       ��o�N�@�            �n@������������������������       �c�VJ/@G             [@                          �:@���U,	@�           ��@������������������������       �	���4�@D           �@������������������������       ��K-�9�@�            �q@                           @˵e�@d           ��@                           @jJT��@V           ��@������������������������       ���I��+@�            0r@������������������������       �u��xޫ@�           ��@                            @u��jc@           �y@������������������������       ��b�Y1@�            �p@������������������������       ��h�;:�@Y            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     t@     ��@      ;@     �L@      |@      X@     Ў@     �l@     P�@     `v@      C@      �?     �W@      a@              0@     @]@      B@     @n@     @Q@      i@      X@      &@             �@@      P@              @      M@      *@     @X@      @@     �R@     �B@      @              2@      C@              @      E@      $@      R@      "@      H@      3@                      "@      ;@                      @@      @      P@      @      @@      0@                      "@      &@              @      $@      @       @      @      0@      @                      .@      :@              �?      0@      @      9@      7@      :@      2@      @              $@      7@                      ,@              5@      ,@      9@      0@      @              @      @              �?       @      @      @      "@      �?       @       @      �?      O@      R@              $@     �M@      7@      b@     �B@     �_@     �M@      @              3@      =@                      6@             �W@      $@      Q@      7@                      "@      @                      1@              "@      @      >@      ,@                      $@      7@                      @             �U@      @      C@      "@              �?     �E@     �E@              $@     �B@      7@      I@      ;@     �M@      B@      @              $@      *@                      &@              (@      �?      :@      @       @      �?     �@@      >@              $@      :@      7@      C@      :@     �@@     �@@      @      $@     @l@     �x@      ;@     �D@     �t@      N@     @�@      d@     �@     `p@      ;@      $@     �c@     @n@      1@      8@     �n@      G@     @n@     �_@     p@     �f@      2@       @      :@      D@               @     �P@      �?      V@      :@      O@     �B@       @       @      5@      9@              �?     �K@      �?      H@      3@     �D@      =@       @              @      .@              �?      &@              D@      @      5@       @               @     �`@     @i@      1@      6@     `f@     �F@     @c@     @Y@     `h@      b@      0@      @     �V@      d@      (@      .@     �b@     �@@      `@     �T@     @d@     �S@      *@       @     �D@     �D@      @      @      ?@      (@      9@      3@     �@@     @P@      @              Q@      c@      $@      1@      V@      ,@     `@     �@@      v@     @T@      "@             �E@     @Z@       @      @      I@      $@     �w@      1@     �o@      G@      @              2@      D@               @      4@      $@     @[@      @     �Q@      *@      @              9@     @P@       @      @      >@             �p@      *@     �f@     �@@       @              9@     �G@       @      (@      C@      @      _@      0@     �X@     �A@      @              4@      C@      @      $@      >@      @     �P@      $@     �P@      0@      @              @      "@       @       @       @      �?     �L@      @     �@@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�6ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�V�\�?@�	           ��@       	                     @�.�+�@e           &�@                          �<@�͝��@b           ��@                           �?
��[(@�           $�@������������������������       ��;u߱@�            @x@������������������������       �^����@           (�@                           �?T�Z �	@h            �d@������������������������       �4i~�~@!            �F@������������������������       �|�P�W�	@G            @^@
                           @�+E���@            �@                           �?%G��c�@�           ��@������������������������       ����γ		@z           Ё@������������������������       �P��p�N@Z            @c@                           @
m�@/             T@������������������������       �R$�(%@#             K@������������������������       ���a��#@             :@                           @7�M��@4           ؚ@                           �?�Y��)@�           (�@                          �4@�E���?�            �v@������������������������       �t��^���?�             n@������������������������       �$c�V�@Q             ^@                           @��A
c@�           �@������������������������       ���o��@�            q@������������������������       �T�ߣb@J           ��@                          �5@��m)�@U           `�@                          �4@>EV��.@�            s@������������������������       �fϴ���@�            @p@������������������������       ��[u	G@            �F@                           �?�G�q��@�            `o@������������������������       ����&�+@D            �Z@������������������������       �L�4�	�@T             b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �q@     8�@      :@      M@     �}@      U@     H�@     `h@     �@     pv@      B@      3@     �i@     �s@      2@     �E@     �t@     �M@      x@     �d@     �x@     �m@      =@      @     �a@     �g@       @      <@     �j@      C@     �m@      Z@     �o@      c@      3@      @     �_@     �e@       @      5@     �g@      8@     �k@     �S@      n@     @^@      *@       @     �F@      J@      �?      @      I@      �?     �X@      $@      X@      ;@       @      @     �T@     �^@      @      2@     �a@      7@      _@      Q@      b@     �W@      &@      �?      .@      .@              @      7@      ,@      *@      :@      .@      ?@      @              @      @                       @      @      @      &@      @      "@              �?      $@       @              @      5@      $@      "@      .@      (@      6@      @      (@     @P@     @_@      $@      .@     �\@      5@     �b@      O@      a@      U@      $@      @     �M@     �Z@      $@      .@     @X@      4@     �a@     �J@     �`@     �S@       @      @     �K@      T@      $@      *@      U@      0@     �V@      E@      Z@      P@       @              @      ;@               @      *@      @      I@      &@      =@      ,@              "@      @      2@                      2@      �?      @      "@      @      @       @      �?      @      0@                      (@      �?      @       @       @      @      �?       @       @       @                      @              @      �?       @              �?             �R@     �m@       @      .@      b@      9@     H�@      =@     P{@     �^@      @             �H@     �c@      @      @      V@      2@     �}@      0@      q@     �P@      @              @     �C@                      .@      @      i@      @      S@      (@                      @      3@                       @             �b@      �?      J@      @                      @      4@                      @      @     �I@       @      8@      @                      E@     �]@      @      @     @R@      &@     Pq@      *@     �h@     �K@      @              5@      M@              �?      4@      &@     @T@      �?      M@      2@      @              5@     �N@      @      @     �J@             �h@      (@     �a@     �B@                      :@     �S@      @       @     �L@      @     `a@      *@     `d@      L@      @              (@     �C@      @       @      8@       @     �X@       @     @W@      4@      @              (@     �@@      @       @      5@             �T@       @     �S@      3@                              @                      @       @      0@              ,@      �?      @              ,@      D@       @             �@@      @      D@      &@     �Q@      B@                      @      6@                      2@       @      6@      @      7@      *@                      $@      2@       @              .@      @      2@       @     �G@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�(�rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�K��KA@�	           ��@       	                   �5@a\�t�@�           d�@                           �?���\�@�           ��@                          �3@�_у��@           �x@������������������������       ���W��@�            �l@������������������������       �ƿç��@b            �d@                          �1@.�8G?@�            �@������������������������       ��	`��@p            @f@������������������������       �?$����@X           ��@
                           �?�}.	N	@�           �@                           �?�x��	@�            �q@������������������������       ��f=�@�            `m@������������������������       �B��j�@            �F@                          �9@I�a��	@           `�@������������������������       �+��a�@            }@������������������������       �j�u��h
@�            �u@                          �5@r��@"           \�@                           �?���k@�           ��@                          �2@B��5�"�?�            �w@������������������������       �z�=��t�?�            �j@������������������������       ���;��?h            �d@                            @)iN�b�@�           X�@������������������������       �&�,�P�@q           @�@������������������������       �)K �@>            �X@                          �<@�-6�%@}           ��@                          �7@��G|9v@G           H�@������������������������       ��)2�v@�            �j@������������������������       �W��Bc@�            Ps@                           @�)��~�@6            �Y@������������������������       �oX���@             C@������������������������       �g�V�@#            @P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@      @@      I@     @~@     �O@     �@     `n@     ��@     `t@      ?@      2@     �k@     Pu@      2@     �B@     �u@     �K@      y@      i@     �u@     �k@      9@       @     �T@     `e@      @      (@     @d@      3@     `p@     �Y@      j@      W@      &@      @      <@     @R@      @      �?     �L@      $@      W@     �E@     �F@     �A@       @      @      0@      B@      �?              9@      @      O@      :@      ;@      <@              �?      (@     �B@       @      �?      @@      @      >@      1@      2@      @       @      @      K@     �X@       @      &@     @Z@      "@     @e@     �M@     `d@     �L@      "@              ,@      <@                      4@              N@      "@     �B@      $@              @      D@     �Q@       @      &@     @U@      "@     �[@      I@     �_@     �G@      "@      $@     �a@     @e@      *@      9@     �f@      B@     @a@     �X@      a@      `@      ,@              E@      @@              @     �I@       @      H@      ,@     �H@      B@      @             �C@      ?@              @      G@      �?      ;@      *@     �C@     �@@      @              @      �?                      @      �?      5@      �?      $@      @              $@     �X@     @a@      *@      6@     ``@      A@     �V@      U@      V@      W@      &@      @      J@     �W@      @      (@     �S@      @     �M@     �E@      M@     �G@      @      @     �G@      F@      @      $@     �J@      ;@      ?@     �D@      >@     �F@       @             �W@     `k@      ,@      *@     �a@       @     h�@     �E@     `z@     �Z@      @              B@     @a@      @       @     �N@      @     |@      0@     �q@     �L@      @              @      E@              @      1@              k@      @     @T@      @      @              @      0@                      &@              a@      @      A@      @      @              @      :@              @      @              T@      �?     �G@                              >@      X@      @      @      F@      @      m@      &@      i@      I@      �?              6@     �V@      @      @      C@      @     `g@      $@      f@      G@      �?               @      @       @              @      �?      G@      �?      9@      @                     �M@     @T@       @      @     �S@       @     �e@      ;@     �a@     �H@       @             �D@      Q@      @      @     �L@       @      d@      9@      ^@     �B@       @              3@     �B@      @              6@      �?     �R@       @     �B@      .@                      6@      ?@              @     �A@      �?     �U@      7@     �T@      6@       @              2@      *@      @       @      6@              &@       @      4@      (@                              @      @       @       @              @       @      &@      @                      2@      @                      4@              @              "@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJo�[*hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��XJ@�	           ��@       	                    �?��b��@y           �@                           �?C����H	@�           ��@                          �<@;Rw@�l@(           �}@������������������������       ���_"��@           Pz@������������������������       ��å�#@!            �L@                          �9@�>{���	@�           �@������������������������       �"��RD	@	           �@������������������������       �y�Rf��
@�            `r@
                           �?�ɛ��@~           p�@                           �?�.��ה@q            `d@������������������������       �,­�@�@7            �S@������������������������       ��K �F@:            @U@                          �2@oaP�o�@           �z@������������������������       �X��Q_�@K            �]@������������������������       ����d�@�            Ps@                           �?��_�l@A           X�@                          �4@���Lu@r           ��@                            �?��Q� @�            0v@������������������������       �'v�Z�?:            �W@������������������������       �^x^@�            @p@                            @փ���@�            �m@������������������������       ��<^K?@�            �i@������������������������       �|����?             @@                          �7@��X̼�@�           �@                          �6@p/�x3@           ��@������������������������       ��&���@�           ��@������������������������       ��US�`@5            @X@                           �?��Yf@�            �r@������������������������       ��� �KI@O            ``@������������������������       �g�Lr~�@f            `e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     @s@     ��@      <@      Q@     �{@      R@     ��@     �i@     ��@     Pv@      B@      ,@     @j@     Pt@      6@      I@     �q@      J@     x@     �d@     x@     �m@      >@      ,@      f@      n@      3@     �C@     `j@      G@      n@     �]@     �p@      f@      <@              G@      R@      �?      &@      M@      �?     �[@      8@     �[@      E@       @              B@     �Q@      �?      @      I@      �?     @[@      6@     @Y@      8@       @              $@       @              @       @               @       @      "@      2@              ,@     ``@      e@      2@      <@      c@     �F@      `@     �W@     @c@     �`@      :@      @     @W@     @a@       @      4@     @^@      3@     �Z@     �O@     �^@     �T@      4@      @      C@      >@      $@       @      @@      :@      7@      ?@      ?@      J@      @             �@@     @U@      @      &@     �R@      @      b@      H@     @^@     �N@       @               @      $@              @      3@             @P@      @     �F@      $@                      @       @              @      &@             �B@       @      0@      @                      @       @                       @              <@      �?      =@      @                      9@     �R@      @       @      L@      @      T@     �F@      S@     �I@       @              @      *@               @      1@             �F@      .@      (@      "@                      4@      O@      @      @     �C@      @     �A@      >@      P@      E@       @      �?     �X@     @o@      @      2@     �c@      4@     �@     �C@     �x@     �]@      @              2@     �U@              @      ;@      @     �q@      *@     @`@      7@      �?              &@      F@              @      *@             `h@       @     �P@      *@      �?                      &@                                      O@              .@      @                      &@     �@@              @      *@             �`@       @      J@      @      �?              @      E@                      ,@      @     @V@      @     �O@      $@                      @     �D@                      (@      @      P@      @      N@      $@                      �?      �?                       @              9@              @                      �?      T@     �d@      @      .@     @`@      *@     v@      :@     �p@      X@      @             �I@     �`@      @       @      R@       @     �r@      $@     �i@      L@      @              E@     @Z@      @      @     �P@      @     �q@      "@     �g@      H@      @              "@      >@              @      @       @      3@      �?      2@       @              �?      =@      =@              @      M@      @      J@      0@     �O@      D@       @      �?      *@      4@              @      =@              ,@      @      ;@      ,@       @              0@      "@              @      =@      @      C@      "@      B@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ;�W@hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?5MBkf@�	           ��@       	                   �<@1�hfn	@�           ��@                           �?�f��3	@�           x�@                           �?	�W���@           �{@������������������������       ��!^�@k             d@������������������������       ���R�`@�            �q@                           @d{b^��	@g           (�@������������������������       �	W�9�Z	@           �{@������������������������       ���2�	@T           h�@
                          �A@�tŶ@y            `i@                            @X�2B{@r             h@������������������������       ���	@;            �[@������������������������       �=�I��@7            �T@������������������������       �������?             $@                          �2@V>[�_�@�           ��@                           �?@���I@�           X�@                           @փc����?�            `q@������������������������       ���:3�v�?x            �f@������������������������       ��>f�*@=             X@                           �?��Ct�@           Py@������������������������       �VQ`�@{            �g@������������������������       ��G#� @�             k@                           �?��r��@�           Ԙ@                           @ݐ:,�@�           x�@������������������������       ��Xh�L�@           0z@������������������������       ���­�@�            �v@                           @��C���@�           0�@������������������������       �޵�`Ӎ@�           P�@������������������������       ��
�L@             <@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        6@     r@     H�@     �B@      H@     �{@     �V@     ��@     �l@     �@     @v@     �@@      5@     `d@     �m@      :@      :@     @n@      M@     `k@     �a@     �p@     �j@      :@      .@     `a@     �j@      8@      5@     @l@      E@     �j@     �]@     `n@     @c@      :@             �K@     @R@      @       @      N@      �?      V@      8@     @X@      @@      @              ,@      :@                      1@             �E@      �?     �F@      *@       @             �D@     �G@      @       @     �E@      �?     �F@      7@      J@      3@       @      .@      U@     �a@      3@      3@     �d@     �D@     �_@     �W@     @b@     �^@      6@       @     �C@      M@      (@       @     �U@      5@      O@      4@     @P@     �L@      @      @     �F@      U@      @      &@      T@      4@      P@     �R@     @T@     @P@      2@      @      8@      8@       @      @      0@      0@      @      6@      7@      N@              �?      8@      5@       @      @      0@      0@      @      5@      7@     �M@                      (@      @              �?      @      &@      @      0@      *@     �E@              �?      (@      .@       @      @      $@      @       @      @      $@      0@              @              @                                              �?              �?              �?     �_@     �s@      &@      6@     �h@      @@     �@     �U@     ��@     �a@      @              9@     �S@      �?      �?     �@@             t@      .@     �d@      E@      �?              *@      ?@                      (@             �a@      �?      Q@      $@      �?              @      1@                      @             �Z@              E@      "@                       @      ,@                      "@              B@      �?      :@      �?      �?              (@     �G@      �?      �?      5@             `f@      ,@     �X@      @@                      @      5@      �?              1@             @Q@      $@      G@      2@                      @      :@              �?      @             �[@      @      J@      ,@              �?     @Y@     �m@      $@      5@     �d@      @@     �}@      R@     w@      Y@      @      �?      J@      ^@      @      (@     �W@      "@      k@      =@     �g@      I@      @      �?      C@     @R@              @     �M@      @     �U@      6@      W@     �A@      @              ,@     �G@      @       @      B@      @      `@      @     �X@      .@                     �H@      ]@      @      "@     �Q@      7@     @p@     �E@     @f@      I@       @              E@      \@      @      "@     �P@      6@      p@      B@     @f@     �H@       @              @      @      �?              @      �?      @      @              �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJa�|rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @-�	˫Y@�	           ��@       	                    �?QI��@u           :�@                          �2@	SA6�@�           ��@                           �?5�O��@x            �f@������������������������       ��0�B@4             S@������������������������       �p�(��@D            @Z@                           �?�{L��B@4           �}@������������������������       ��[LB@�            �u@������������������������       �u�Se-�@R            �`@
                           �?��Aa�	@�           (�@                           �?$.]!�@Q            `a@������������������������       �=��,@             >@������������������������       �b��C��@B            @[@                           �?���2r	@x           ��@������������������������       �$��`��	@�           ��@������������������������       �E}�f˰@�            �x@                          �5@�?i�@=           ��@                            @c:��@�           �@                           �?|>gx2@D           ��@������������������������       ��@b����?�            0u@������������������������       � �3�#@y           �@                          �4@�$� $��?k            �e@������������������������       ��嘌���?^            `c@������������������������       ��6,؊� @             4@                          �<@��7��@�           @�@                           �?X�kzI@W           ؀@������������������������       �>��,�@�            �p@������������������������       ����<@�            �p@                           @5�̈́��@7            @S@������������������������       �K2�5�n@&            �K@������������������������       ��ڇ+��@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@      �@      >@      K@     pz@     @U@     ��@     `k@     ��@     `w@     �@@      .@      l@     �u@      7@     �F@     �q@      P@     pu@      g@     `w@     �p@      =@             @Q@     @Z@               @     �S@      @     `a@      D@      b@     @P@      @              @      3@               @      6@              O@      @     �G@      2@                       @      $@                      ,@              =@      @      &@      @                      @      "@               @       @             �@@       @      B@      &@                     �O@     �U@              @      L@      @     @S@     �A@     �X@     �G@      @              G@      R@              @     �F@       @      E@      =@     �N@      D@      @              1@      ,@               @      &@       @     �A@      @     �B@      @       @      .@     �c@     �n@      7@     �B@      j@      N@     �i@      b@     �l@     @i@      7@      @      2@      (@              @      :@      @       @      ;@      4@      1@      @               @      �?                      "@       @              @      @      @              @      0@      &@              @      1@      @       @      7@      ,@      &@      @      (@     @a@      m@      7@      ?@     �f@     �K@     @i@     @]@      j@      g@      4@      (@     �Z@     @d@      6@      8@     @`@      F@      ^@      V@     �a@      b@      1@              @@     �Q@      �?      @      J@      &@     �T@      =@      Q@      D@      @       @     �R@     @l@      @      "@      a@      5@     ��@     �A@     �{@     �Z@      @              D@     �`@              @     �N@      $@     �}@      0@     pr@      K@      @              @@     �_@              @      I@      $@     �x@      .@     �l@      H@       @              @     �E@              @      *@      �?     �g@      @      P@      &@      �?              :@      U@               @     �B@      "@     �i@      "@     �d@     �B@      �?               @      @                      &@              S@      �?      P@      @       @               @      @                      @             @Q@      �?     �M@      @                                                      @              @              @      �?       @       @     �A@      W@      @      @      S@      &@     �d@      3@     �b@     �J@               @      8@      U@      @       @      K@      &@     �c@      1@     `a@     �D@               @      1@      H@      �?              ;@      �?     @S@      $@     �O@      7@                      @      B@      @       @      ;@      $@     �T@      @      S@      2@                      &@       @      �?      �?      6@               @       @      (@      (@                      @       @              �?      3@              @      �?      "@       @                       @              �?              @               @      �?      @      @        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ6SShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?곈�]Q@�	           ��@       	                   �3@�*���@:            �@                           @K���r�@�           ��@                           �?׀�W�@�            �o@������������������������       ���yX-�@<             X@������������������������       �q/��E@b            �c@                           @]��rK @�            �y@������������������������       ����Y�V�?�            �s@������������������������       �g�wо@B             X@
                           �?�I���*@�           ̐@                           �?e���_�@�            �w@������������������������       �|a���9@^            `c@������������������������       �o�ʌ��@�            @l@                           @�I�y��@�           ��@������������������������       �d���v	@�            �v@������������������������       �H�e�]@�            �t@                          �:@��ז�|@Z           �@                            @ؐ�z��@v           ��@                          �9@�C�|��@1           ��@������������������������       �Xr�|�v@           l�@������������������������       ����@�"@*            �Q@                           �?�����@E           �@������������������������       �<�S�"@S            �a@������������������������       ��m�>�c@�            Pw@                            �?�)�L&	@�            �u@                           �?���$�@A            @Z@������������������������       �|%��b�?             "@������������������������       ��9���@:             X@                            @�_FJ�@�            �n@������������������������       ��Dɯ}�@]            �a@������������������������       ��붜@F             Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     x�@      <@     �I@     �z@     �W@     ��@      j@     H�@      x@      @@       @     �Y@     �o@      *@      :@     �h@      C@     �@     �U@     ps@      g@      &@      @      4@      U@      �?      @      H@      @      r@     �@@     �Z@      P@      @      @      (@     �A@                      5@      @      Q@      <@      B@     �D@      @              @      &@                      @      @      B@      $@      1@      @              @      @      8@                      .@       @      @@      2@      3@      A@      @               @     �H@      �?      @      ;@             �k@      @     �Q@      7@                       @      C@      �?              0@              g@      @      I@      0@                      @      &@              @      &@             �B@      �?      4@      @              @     �T@     `e@      (@      7@     �b@      @@     �j@      K@     �i@      ^@       @      �?      =@     �I@              "@      E@      @     �\@      0@     @T@      A@              �?      2@      (@              @      4@      �?      3@      *@      D@      9@                      &@     �C@              @      6@       @      X@      @     �D@      "@              @      K@      ^@      (@      ,@     �Z@      =@     �X@      C@      _@     �U@       @      @     �C@     @S@      $@       @     �J@      7@      8@      =@     �C@      L@      @              .@     �E@       @      @     �J@      @     �R@      "@     @U@      >@      @      *@      g@      s@      .@      9@     �l@     �L@     �@     @^@      @      i@      5@      @     �a@      q@      (@      .@     �e@      E@     `}@     �W@     �{@      a@      3@      @      [@     �f@      (@       @     @Z@     �@@     `u@     �P@     �u@     �V@      1@      @     @Y@     �d@      (@       @      Z@      6@     u@      N@      t@     �V@      1@              @      0@                      �?      &@      @      @      7@      �?              @      A@      W@              @      Q@      "@      `@      <@      X@      G@       @              &@      @@               @      @              J@      @      :@      "@              @      7@      N@              @      P@      "@      S@      8@     �Q@     �B@       @      @      E@      >@      @      $@      M@      .@      C@      ;@     �L@     �O@       @              @      @       @              9@      "@      *@      &@      4@      *@      �?                       @                      �?               @              @                              @      @       @              8@      "@      &@      &@      0@      *@      �?      @      B@      9@      �?      $@     �@@      @      9@      0@     �B@      I@      �?      @      2@      *@              @      :@      @       @      @      =@      <@              @      2@      (@      �?      @      @      �?      1@      &@       @      6@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJG�LchG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @j�)��N@�	           ��@       	                    �?1��p��@�           V�@                           �?"��*��@�           D�@                           �?T�yh!�@6            @������������������������       �"MӠ��@|            `h@������������������������       �y�#�`@�            �r@                            �?��դCt	@�           ��@������������������������       �7<4v��@�            Ps@������������������������       ��X��Z	@�           `�@
                           �?B�o��@�           Ђ@                          �<@�S�AU�@n            �e@������������������������       ���U��@g            �c@������������������������       ��1P�E�?             *@                           �?�uN�2)@           �z@������������������������       ��&�Y@             @@������������������������       ���@�h�@	           �x@                           �?�N0�@)           x�@                          �4@tRM��� @k           @�@                            @۸�"���?�            `u@������������������������       �m:V���?�             r@������������������������       ��h�ܻ�?%             K@                            �?����1@�            @j@������������������������       ���xQ@             B@������������������������       �Ѓ�Y@s            �e@                            �?_mB@�           ؑ@                          �1@'hٔ$1@�           ȃ@������������������������       �
_���?M            @^@������������������������       ��^_���@4            �@                           �?Bh��@=           �@������������������������       ���qY@�             n@������������������������       ��㸆�C@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        "@     �t@     ��@      @@     �M@      }@      U@      �@     �j@     `�@     0u@      <@       @     `n@     �t@      9@     �D@     0u@      O@     @w@      g@     v@     �m@      5@       @      g@     �o@      7@      >@     �p@      F@     @l@      `@     �n@      g@      4@              O@     @U@       @      @     �P@      �?     @Y@      :@      W@     �I@      @              7@      ;@                      6@              L@      @      G@      ,@      @             �C@      M@       @      @     �F@      �?     �F@      6@      G@     �B@      �?       @     �^@     �d@      5@      9@     `i@     �E@     @_@     �Y@     @c@     �`@      0@      �?      G@      7@      @      "@      P@      @     �E@      C@     �D@      ;@      @      @     @S@      b@      0@      0@     `a@     �B@     �T@     @P@     @\@     �Z@      $@              M@     @T@       @      &@     @Q@      2@     @b@     �K@     �Z@      K@      �?              1@      .@              �?      7@      @      Q@      @     �@@      @                      0@      ,@              �?      1@      @     �P@      �?     �@@      @                      �?      �?                      @              �?      @                                     �D@     �P@       @      $@      G@      *@     �S@      I@     �R@     �H@      �?              @      @              @      �?      �?      �?      @      @      @                     �B@      O@       @      @     �F@      (@     @S@     �F@     �Q@     �E@      �?      �?     �V@     �m@      @      2@     �_@      6@     ��@      >@     �z@     @Y@      @              (@     �R@       @       @      >@      @     �p@      @     `a@      2@      �?              @     �C@               @      (@             @h@      @     �S@      @      �?              @      C@              �?      "@              d@      @      Q@      @      �?              �?      �?              �?      @              A@              &@      @                      @     �A@       @              2@      @     �Q@       @      N@      (@                              @       @              @       @      *@              @      @                      @      >@                      (@       @      M@       @     �K@      "@              �?     �S@     �d@      @      0@     @X@      2@     pv@      9@      r@     �T@      @             �I@      Y@      �?      $@     �D@      $@     �f@      0@      e@      K@      �?                      .@              @      @              L@             �A@      @                     �I@     @U@      �?      @     �A@      $@     @_@      0@     �`@     �H@      �?      �?      <@     @P@      @      @      L@       @     @f@      "@      ^@      =@      @      �?      &@      8@      @      @      @@      �?      T@      @      L@      5@      @              1@     �D@      �?      @      8@      @     �X@      @      P@       @       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�5=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Py��+G@�	           ��@       	                    �?	�B�@           ��@                          �2@�`rW\}@0           @}@                           �?���N�@M             \@������������������������       ��筱:� @&             M@������������������������       ��'�*��@'             K@                          �<@�v4* @�            @v@������������������������       �}��(�@�            �r@������������������������       �>o�y�@"            �J@
                           @Q�g��@�           ؈@                            �?O��ހ$@f           X�@������������������������       �A�[K���?]             d@������������������������       ��$oQJ�@	           �z@                          �:@�7��@�             j@������������������������       ����^z9@u            @g@������������������������       ��~~�x @             6@                          �1@�b��vO@�           ��@                           @� �~��@�            �u@                           �?��C��@j            `f@������������������������       �ӯ�jI�@+            �U@������������������������       ��Q��V�@?            @W@                           �?����?p            @e@������������������������       �=���^ @;            �W@������������������������       �*�����?5             S@                           @�r���@�           ��@                           @-�lBw@           ��@������������������������       ��V����	@�           ��@������������������������       ����I�F@           �@                           @���",	@�            �q@������������������������       ����o�S	@y            �g@������������������������       �&tu�(@9            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �r@     H�@     �B@      K@      {@     �S@     ��@     @l@     ��@     pu@      8@      �?     �T@     �e@              &@     �X@      &@     �}@      E@     @r@     @R@      @      �?      H@     �P@              @      H@       @     �[@      A@     �Z@     �E@       @              @      5@                      .@             �D@       @      8@      @                      �?      *@                      @              7@      �?      *@                               @       @                       @              2@      �?      &@      @              �?     �F@      G@              @     �@@       @     @Q@      @@     �T@     �B@       @      �?      A@     �C@              @      <@       @     �P@      ;@      S@      7@       @              &@      @               @      @               @      @      @      ,@                     �A@      [@              @     �I@      "@     �v@       @      g@      >@       @              =@     @R@                     �D@       @      r@       @     �^@      7@      �?                      =@                      @      @      V@              ;@      @      �?              =@      F@                     �A@      @      i@       @     �W@      1@                      @     �A@              @      $@      �?     �R@      @     �O@      @      �?              @      ?@              @      $@             @R@      @      J@      @      �?                      @                              �?      �?      @      &@       @              7@     �j@     �w@     �B@     �E@     �t@     �P@     ��@      g@     ��@     �p@      4@              3@      I@      �?       @      7@             �`@      4@     @S@      8@                      ,@      ;@      �?      �?      0@             �H@      3@     �@@      3@                      @      $@      �?              $@              8@      .@      "@      *@                      $@      1@              �?      @              9@      @      8@      @                      @      7@              �?      @              U@      �?      F@      @                      @      1@              �?      @              I@      �?      *@      @                      �?      @                      @              A@              ?@      �?              7@     �h@     �t@      B@     �D@     �s@     �P@     �y@     �d@     �|@     �n@      4@      0@     �d@     Pr@     �A@     �D@     q@      L@     @w@     �^@     �y@     `k@      &@      0@     @\@     �d@      >@      ?@     �h@     �E@     �`@      Z@     �h@     @b@      $@              K@     �_@      @      $@      S@      *@      n@      2@      k@     @R@      �?      @      =@     �A@      �?             �C@      &@     �B@      E@      G@      ;@      "@      @      5@      ;@      �?              ;@      $@      0@      B@      2@      4@      @               @       @                      (@      �?      5@      @      <@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��:9@�	           ��@       	                    �?+R�qh�@�           z�@                            �?w�\{ @�            �@                          �8@A��7+@�            �m@������������������������       ��; ]��@m            @e@������������������������       ��#����@$            �P@                           �?���@1           @}@������������������������       �ƿ�K@�            `u@������������������������       ���(�l@M            �_@
                          �4@W�CT�	@�           ��@                           @ ieo>@y           ��@������������������������       �P�3�P�@k            �@������������������������       ����@             7@                           �?}Pط��	@W           0�@������������������������       ���cU}@�            Pp@������������������������       ���:.�	@�           �@                          �4@�����@6           0�@                           @�N�@8           x�@                            �?���i>@            `h@������������������������       ��5�K�@L            @]@������������������������       ����k�@3            �S@                           �?0A���1@�           `�@������������������������       ���3���?�            @o@������������������������       �r+[�L@            {@                           @�z���@�           �@                            @�`a]@D           P@������������������������       �Y���@           �y@������������������������       ��{��y��?1            @V@                            �?��;l�5@�            �r@������������������������       �&
��@,            �P@������������������������       ��� �L@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     `q@      �@      ;@     �O@     p{@      R@      �@     �k@     @�@     �u@      ;@      7@     �h@     `u@      4@     �J@     �r@     �L@      y@      g@     y@     �m@      4@      �?     �P@     �Z@       @      @     �Q@      @     �e@      B@     `e@     �P@       @      �?      8@     �C@              �?      7@      �?      J@      @      R@      ,@       @              (@      8@              �?      6@      �?      H@      @     �J@      @              �?      (@      .@                      �?              @       @      3@      $@       @             �E@     �P@       @      @      H@      @     @^@      =@     �X@     �J@                      >@      K@       @      @     �A@              T@      :@     �P@     �F@                      *@      *@                      *@      @     �D@      @      @@       @              6@     �`@     �m@      2@     �H@      l@     �J@     �l@     �b@     �l@     �e@      2@      "@      B@     @Q@      @      &@     �T@      &@     �]@      G@     �_@      G@      @      @      A@     �P@      @      &@     @S@      "@     �\@     �F@     @_@      G@      @      @       @       @                      @       @      @      �?      �?              @      *@      X@     �d@      &@      C@     �a@      E@     �[@     �Y@      Z@     �_@      (@       @      &@     �C@      �?      0@      D@      @     �D@      4@      >@     �J@      @      &@     @U@      `@      $@      6@     �Y@     �B@     �Q@     �T@     �R@     @R@      "@             �S@     �m@      @      $@     �a@      .@     p�@      C@     p{@     �[@      @              @@     �_@      �?      @     �B@      @     @x@      "@     �k@      M@      �?              (@     �A@                      $@      @     @S@             �G@      &@                      @      6@                      @             �H@              ;@      "@                      @      *@                      @      @      <@              4@       @                      4@     �V@      �?      @      ;@             ps@      "@     �e@     �G@      �?              @     �@@                      @             `a@       @      L@      $@      �?              ,@      M@      �?      @      8@             �e@      @     �]@     �B@                     �G@      \@      @      @     �Z@      (@     @i@      =@     @k@      J@      @              A@     �J@      �?       @     �P@       @     �b@      ,@     `b@      :@      @             �@@     �I@      �?       @      J@      �?     �[@      ,@     @]@      9@      @              �?       @                      ,@      �?      D@              >@      �?                      *@     �M@      @      @      D@      $@     �I@      .@     �Q@      :@      �?              @      @      @              @      @      1@      @      (@      @                      @     �J@       @      @      A@      @      A@      $@     �M@      5@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�e�ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?W�#�:@�	           ��@       	                    �?Y��8��@           ��@                           �?2�	��@�            �@                          �:@�����@�            �l@������������������������       ���5�@t            `f@������������������������       ����[�@            �H@                           @�w��@           �y@������������������������       �����@l            �d@������������������������       ���܇ @�            �n@
                           �?ɋ�� @s           ��@                           �?�P!4�@�            �p@������������������������       �%��=��@?             Y@������������������������       ���Xs@e            �d@                           @��� �@�            �v@������������������������       �Q����� @�            �n@������������������������       �b#g�E@J            �^@                          �5@����R'@�           ��@                           �?m�	��@u           `�@                           �?�cm�0�@A           �~@������������������������       ���- @j            �d@������������������������       ���6�M@�            @t@                          �4@P:�Ly�@4           p�@������������������������       ���&��-@�           ��@������������������������       �� :��:@[             b@                           �?�bG�.	@2           �@                          �6@Q����	@�           �@������������������������       �y���k�@@             [@������������������������       �ׅZ|

@L           P@                          �7@v3��%_@�           ��@������������������������       ��"���p@�            �m@������������������������       ��3��fs@	           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     r@     ��@      <@     �I@     }@      S@     `�@      i@      �@      x@      :@       @     �S@     �e@      @      &@     �[@      *@      |@     �B@     �r@     �W@       @       @      B@     �U@       @       @      M@      @      n@      7@     �^@     �K@               @      3@     �@@       @      @      =@      �?     �E@      0@      E@      B@                      3@      =@       @      @      :@      �?     �B@      *@      A@      .@               @              @               @      @              @      @       @      5@                      1@      K@              @      =@      @     �h@      @     @T@      3@                      (@      4@              �?      0@      @     �R@      �?      8@      .@                      @      A@               @      *@       @     �^@      @     �L@      @                      E@      V@      �?      @      J@      @     @j@      ,@     �e@      D@       @              6@     �D@              @      B@              O@      (@     �P@      7@      �?              $@      (@                      &@              ;@      �?      ?@      @      �?              (@      =@              @      9@             �A@      &@     �A@      0@                      4@     �G@      �?              0@      @     �b@       @     �Z@      1@      �?              1@      >@                      *@      @     @[@             @P@      @                      @      1@      �?              @             �C@       @      E@      ,@      �?      7@     `j@     @x@      9@      D@     0v@     �O@     P�@     `d@     �@     0r@      8@      "@     �Q@      l@      @      4@      d@      8@     pv@     �P@     �r@     �_@      @      "@      E@     �T@      @       @      V@      "@      R@      B@      S@      N@      @      @      0@     �E@      @       @      >@      @      ,@      &@      1@      6@              @      :@     �C@      �?      @      M@      @      M@      9@     �M@      C@      @              =@     �a@      �?      (@      R@      .@     �q@      ?@     �k@     �P@      @              ;@     �^@      �?      $@     �M@      @     �o@      9@     �e@     �N@                       @      3@               @      *@      &@     �A@      @      H@      @      @      ,@     �a@     �d@      3@      4@     `h@     �C@     `h@      X@      j@     �d@      2@      (@      Q@     �T@      ,@      "@     �\@      <@     �J@     �L@     �N@     �W@      1@       @      0@      :@              �?      ,@       @      @      $@      *@      ,@              $@      J@      L@      ,@       @      Y@      4@     �H@     �G@      H@      T@      1@       @      R@     �T@      @      &@     @T@      &@     �a@     �C@     `b@     �Q@      �?              A@      A@       @      @      9@      @     �P@      @      D@      5@               @      C@      H@      @       @      L@      @     �R@     �@@     �Z@      I@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�kS�	Q@�	           ��@       	                   �4@��J���@u           B�@                           �?����L@/           h�@                           @&Y&���@h           0�@������������������������       �����V�@           �z@������������������������       �q��N-	@S            �^@                           �?�]ƿ�Z@�            pt@������������������������       �Ƈ���,@L            @`@������������������������       �%Cq,p�@{            �h@
                           �?+�p'A	@F           Д@                           �?����:r	@�           (�@������������������������       ���v7Q�@�             v@������������������������       ����*��	@�           P�@                           �?�]�ɽ@�            �r@������������������������       �^{d�@6            �S@������������������������       ��෋d"@�            `k@                           �?m�B��$@7           ��@                           @��I�� @b           P�@                          �8@�O;��?�            0u@������������������������       ��F�����?�            �r@������������������������       �>@XBQ�?            �D@                           �?�DiwK�@�            �j@������������������������       �F2rVI:@L            �_@������������������������       ��,��;@7            @V@                          �<@�W �A@�           ��@                           !@�&4.9�@�           ��@������������������������       �:�o�y@�           h�@������������������������       �>�V���?             *@                          �=@�l��@.            �U@������������������������       ��e�M`�?             :@������������������������       �00��E@             �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     ��@      C@     �H@     p~@      T@     ��@      i@     P�@     �v@      <@      6@     �j@     �t@      :@     �A@      u@      N@     �v@      d@     �x@     `n@      :@      @     �I@      ^@      @      $@     �\@      1@     �k@      O@     �f@      T@      &@      @     �B@      P@      @      @     �S@      1@      ^@     �B@      ^@      K@      &@       @      ;@     �F@      @       @     �K@      (@     �Z@      <@      Y@     �F@      �?      �?      $@      3@               @      7@      @      ,@      "@      4@      "@      $@              ,@      L@      �?      @     �B@              Y@      9@      O@      :@                      @      :@      �?              4@             �C@      (@      ,@      &@                      @      >@              @      1@             �N@      *@      H@      .@              3@      d@      j@      4@      9@     �k@     �E@     @b@     �X@     �j@     `d@      .@      3@     �`@     �e@      4@      6@      f@      >@     �Y@     �R@      b@     �_@      *@       @      >@      N@       @      @     �O@       @      K@      <@     �N@     �D@      @      1@     �Y@     @\@      2@      1@     @\@      <@     �H@     �G@      U@     @U@      "@              =@     �A@              @     �F@      *@     �E@      8@     �P@     �B@       @              @      @                      @       @      5@      @      9@      @                      8@      =@              @      C@      &@      6@      2@      E@      >@       @             �V@     �j@      (@      ,@     �b@      4@     p�@     �C@      x@     �^@       @              (@      R@               @      =@       @     0q@       @     @^@      ;@                      @      F@                      *@       @      g@             �Q@      (@                      @     �E@                      (@      @     �d@             �L@      $@                              �?                      �?      @      2@              ,@       @                      @      <@               @      0@             �V@       @      I@      .@                      @      3@               @       @             �N@      �?      9@      @                      �?      "@                       @              =@      @      9@      $@                     �S@     �a@      (@      (@     �^@      (@     �w@      ?@     pp@      X@       @              M@     @a@      "@      "@     �Y@      (@     pw@      ?@     �o@     �R@       @              L@     @a@      "@      "@     �X@      @     pw@      ?@      o@     �R@       @               @                              @      @                      @                              4@      @      @      @      4@              @              &@      5@                      *@       @                      @                              @      @                      @      @      @      @      .@              @               @      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ1�UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@����L@�	           ��@       	                    �?-�/&��@R           �@                           @��+��@�           �@                            �?�St��@�            �u@������������������������       �����@>             Y@������������������������       �Rr>"��@�            �n@                            �?��l�
	@           �x@������������������������       �7c���@L            �]@������������������������       �*�T��	@�            @q@
                           �?p24��P@u           ��@                           �?��b�y�@�           H�@������������������������       �
ÆfBd�?�            �r@������������������������       ��Xwȥ�@           �y@                            �?s5�~��@�           ��@������������������������       �
ة��� @z            `j@������������������������       ����1@C           (�@                           @�9I��@H           �@                          �9@{���o	@�           h�@                            �?��s�:�@�           �@������������������������       �����@t            �f@������������������������       �ϸ$"]@           �z@                           �?N�����	@C           �@������������������������       �8U	A�	@�            Py@������������������������       ����q�@D             Z@                           �?���x��@�           X�@                           �?�Ρ�x@q            �e@������������������������       ��(_�+@=             X@������������������������       �d��m @4            �S@                           @�����\@           �{@������������������������       ��W;@           �z@������������������������       �Nɱ���@             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      t@     (�@      <@     �K@     �|@     �V@     <�@     @k@     x�@     pv@      <@      @      _@      r@       @      ;@     �k@      C@     ��@     �W@     �}@      e@      $@      @      Q@      Y@      @      0@     �\@      2@     @`@     �J@     ``@      W@       @      @      ?@     �H@      �?       @     �C@      �?     �R@      :@     �S@      B@      @                      (@                      (@              @@      @      ;@      (@      �?      @      ?@     �B@      �?       @      ;@      �?      E@      6@     �I@      8@       @      �?     �B@     �I@      @      ,@     �R@      1@      L@      ;@     �J@      L@      @              3@      (@              �?      8@      @      ,@       @      5@      (@      �?      �?      2@     �C@      @      *@     �I@      $@      E@      3@      @@      F@      @              L@     �g@      @      &@      [@      4@     p�@     �D@     �u@     @S@       @              9@      T@      @      @     �N@       @     @t@      3@     �a@     �F@      �?              *@      ,@              @      .@       @     �g@      @      I@      $@                      (@     �P@      @      �?      G@      @     �`@      ,@     @W@     �A@      �?              ?@      [@      �?      @     �G@      (@     �p@      6@      i@      @@      �?              @     �@@                      @      @     �V@      @      N@       @                      :@     �R@      �?      @     �E@      @     �e@      3@     �a@      8@      �?      (@     �h@     �l@      4@      <@     `m@      J@     �s@      _@     @s@     �g@      2@      $@     `c@     �c@      $@      ;@     @e@      G@     @a@     @Y@     @d@     �^@      0@      �?     @U@      X@       @      0@     �[@      3@     �U@     �G@     �V@     �C@      @      �?      ;@      :@              $@      :@      @      A@      3@      2@      (@      @              M@     �Q@       @      @     @U@      0@      J@      <@      R@      ;@       @      "@     �Q@      N@       @      &@     �M@      ;@      J@      K@      R@      U@      "@      "@      M@      H@       @      &@      F@      8@      @@      F@     �L@     �P@      "@              (@      (@                      .@      @      4@      $@      .@      1@               @     �E@     @R@      $@      �?     @P@      @     �f@      7@     @b@     �P@       @       @       @      3@                      @      @     �O@      @     �I@      1@               @       @      $@                      @              E@       @      8@      @                              "@                      @      @      5@      @      ;@      (@                     �A@      K@      $@      �?      M@      @     �]@      2@     �W@      I@       @             �@@     �J@      @      �?     �K@       @      ]@      0@     �W@      I@       @               @      �?      @              @      �?       @       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ4�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�����A@�	           ��@       	                    @!v�G@�           �@                            �?�BfĐe@G           ��@                           �?�s��<�@�            �p@������������������������       ��t:�[@3            �S@������������������������       �4(&
�_@~            �g@                           �?d,K�@�           p�@������������������������       �a���@~            @j@������������������������       ���HB��@           �{@
                           �?�7? �@E           P�@                          �1@�r�5��?�            �t@������������������������       ���q����?`             b@������������������������       �)�xF���?�            @g@                           @��t�W�@d           ��@������������������������       �����5@Q            �a@������������������������       �r�,��@            y@                           @fg�`@F           ��@                           �?�P�n<	@F           ��@                           @����X	@�           �@������������������������       �I؟	@O           ��@������������������������       �(
��@?            @Z@                           �?�8����@�            �q@������������������������       �����X6@R            �_@������������������������       �O�ɇ�@f            �c@                          �7@�ul�@            �@                          �5@OQ�CCo@�            �v@������������������������       �g�9�@b             b@������������������������       ���ȷ�!@�            �k@                           �?X:��@            {@������������������������       ��4�f;@O            @_@������������������������       �������@�            Ps@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      q@     �@      ;@     �L@     �@     �U@     Џ@     �k@     0�@     �u@      =@       @     �W@     �k@      $@      5@     �g@      7@     ��@     �P@     �w@     �`@      @       @     �J@      `@      "@      ,@      a@      2@      l@     �H@      h@     �U@      @              ,@      F@              �?     �C@      @     �Q@      (@     �O@      2@      @               @       @                      (@       @      ?@      @      1@      @                      (@      B@              �?      ;@      @     �C@       @      G@      .@      @       @     �C@      U@      "@      *@     @X@      *@     @c@     �B@      `@     @Q@       @              0@      *@               @      ;@      �?      S@       @     �I@      0@               @      7@     �Q@      "@      &@     �Q@      (@     �S@      =@     �S@     �J@       @             �D@     �W@      �?      @      K@      @     �y@      2@     �g@     �G@                      "@      @@               @      (@             @h@      @     �P@      &@                      @      (@               @      @              U@      �?      ?@      @                      @      4@                      @             �[@      @      B@      @                      @@     �O@      �?      @      E@      @     �k@      ,@      _@      B@                      ,@      :@                      @      @      J@      @      ;@      @                      2@     �B@      �?      @     �A@              e@       @     @X@      >@              &@     �f@      r@      1@      B@     @t@     �O@     �w@     `c@     pz@     �j@      7@      $@     �`@      f@      $@      <@      l@      J@     @d@      `@      j@      d@      4@      $@     �\@     �a@      $@      9@     �e@      @@     �Y@     �Z@     �d@     �`@      2@      @      Z@      `@      "@      9@     @c@      ;@      W@     @T@     �d@     @_@      &@      @      $@      ,@      �?              2@      @      $@      9@      �?      $@      @              5@      A@              @      J@      4@      N@      7@     �E@      9@       @               @      &@               @      9@      @      @@      (@      3@      &@      �?              *@      7@              �?      ;@      .@      <@      &@      8@      ,@      �?      �?     �F@     �\@      @       @      Y@      &@      k@      :@     �j@      K@      @              4@     �Q@      @      �?     �F@      @      ]@      @     @U@      ,@      @              @      A@              �?      &@      @      E@       @      D@      @      @              1@      B@      @              A@       @     �R@      �?     �F@      $@              �?      9@      F@      @      @     �K@      @     @Y@      7@     @`@      D@                      @      0@                      @       @      E@      @     �H@       @              �?      6@      <@      @      @      I@      @     �M@      1@     @T@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ\�C\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?<�"\@�	           ��@       	                    �?t��2D	@           ��@                          �;@V����@4           �~@                           �?�CVj��@            z@������������������������       �Z���@z             i@������������������������       ������@�            �j@                            �?�zg�X@)            @R@������������������������       ����w&�@            �C@������������������������       �BD�Q�D@             A@
                           �?���=e�	@�           �@                            �?N�b�n�@           �y@������������������������       ����%�@E            @\@������������������������       �_��'pi@�            �r@                           �?�y�7�	@�           0�@������������������������       �It$�H	@�            �m@������������������������       �����	@8           �@                           @F�S�@�           ��@                          �9@�6�a6�@           `�@                           �?����w'@8           �}@������������������������       �	i)�@�            @i@������������������������       �xCNj@�             q@                           �?���gF@G             \@������������������������       �NC��2x@             E@������������������������       �4�o��@,            �Q@                            �?��v"�@?           <�@                           �?\A3��@�            �v@������������������������       ��ٝ��N�?O            �_@������������������������       ���x؇"@�            @m@                          �4@�n*F�@P           ��@������������������������       �@����G@�           x�@������������������������       ��^��|m@w           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �s@     8�@      @@     @P@     �|@     �S@     `�@     `m@      �@     �t@      7@      1@     `e@     Pq@      :@     �E@     �n@      I@      l@     �a@     `o@     �f@      ,@      @     �I@      X@      @      &@     @P@       @      V@      @@     @V@     �G@       @              F@      S@      @      @      O@              U@      <@     �S@      ?@       @              2@      ;@      @      @     �@@              H@      2@     �A@      ,@                      :@     �H@               @      =@              B@      $@      F@      1@       @      @      @      4@              @      @       @      @      @      $@      0@              @       @      $@               @      @       @                       @      .@                      @      $@               @                      @      @       @      �?              ,@      ^@     �f@      7@      @@     �f@      H@      a@     �[@     @d@      a@      (@      @      7@      R@      @      .@     �Q@      (@      R@      B@      K@     �I@      @              $@      0@              @      4@      @      <@      ,@      @      @      �?      @      *@      L@      @      &@      I@      @      F@      6@     �G@     �F@       @      &@     @X@     @[@      3@      1@     �[@      B@     @P@     �R@      [@     @U@      "@      @      A@      G@      "@      �?      ;@      *@      3@      :@      5@     �B@       @       @     �O@     �O@      $@      0@      U@      7@      G@     �H@     �U@      H@      @             �a@      s@      @      6@     `j@      <@     X�@      W@     H�@     �b@      "@             �H@     �T@      �?      $@     �P@      $@     �b@     �H@     @]@     �I@      @              A@     �Q@      �?       @      I@      @     �a@      @@     �X@      A@      �?              *@      =@      �?      @      ;@      @     �I@      1@     �E@      *@      �?              5@     �D@              @      7@      @     �V@      .@     �K@      5@                      .@      (@               @      0@      @      "@      1@      3@      1@       @              @      @                      @      �?       @      �?      @      ,@                       @      "@               @      "@       @      @      0@      (@      @       @             �W@      l@      @      (@      b@      2@     ��@     �E@     @y@     �X@      @              9@     �G@       @      �?      8@      @      c@      *@     �O@      ?@                              "@      �?              @       @     �R@      @      8@      @                      9@      C@      �?      �?      3@      �?     @S@      "@     �C@      8@                     @Q@      f@      @      &@     @^@      .@     �}@      >@     Pu@      Q@      @              @@     �W@       @      @      G@      �?     @s@      0@     �f@      =@       @             �B@     �T@      �?      @     �R@      ,@      e@      ,@     �c@     �C@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @[���a�@�	           ��@       	                    �?u�:��_@�           ��@                          �6@�#D@G           ��@                           �?�ۼ
�5@�           ��@������������������������       ����*@�            `u@������������������������       ��Fq��J@�            �q@                           �?���n(�@�            �r@������������������������       �B�R�j@U            @a@������������������������       �Xvn�a>@a            @d@
                           @G�d}/6@�           �@                          �4@��0�@0           X�@������������������������       ��Ě�k@�            �w@������������������������       ���:NO.	@P           ��@                           @
�9ڈo@W           p�@������������������������       ��a�M�@H           ��@������������������������       ���<��@             9@                          �3@J[=Y9@�           Б@                           �?;�uT�@�            0y@                           �?Q�O�a�@�            �i@������������������������       �"�\�@5            @U@������������������������       �$zU�C@M            @^@                          �1@���ʆ@y            �h@������������������������       ����eI @6             U@������������������������       �5��{�a@C            @\@                          �<@��W���@�           �@                          �:@ar�?7�@�           h�@������������������������       �ܦ�0�@c            �@������������������������       ��F+&`�@2            @S@                           �?v�}���@M             ]@������������������������       ��c?���@             8@������������������������       ��d_Ih�@=             W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     p�@      =@      I@     �z@     �P@     ,�@     �i@     h�@     pv@      4@      @     �g@      z@      .@      ;@     �r@      I@     ��@     @a@     H�@     �n@      &@      �?     �F@     @b@      @      @     �Q@      (@     �t@      9@     �j@     �P@                      6@     �W@      �?      �?     �D@      @     �p@      .@     �b@      ;@                       @      H@      �?      �?      @@      @     �d@      (@     �M@      &@                      ,@      G@                      "@              Z@      @     �V@      0@              �?      7@      J@      @      @      >@      @     �P@      $@     @P@      D@              �?      2@      ?@              @      1@              ,@      @      ;@      8@                      @      5@      @              *@      @     �J@      @      C@      0@              @     @b@      q@      &@      7@     `l@      C@     �z@     @\@     0y@      f@      &@      @     @X@      a@       @      (@      a@      =@     �]@     @V@     @c@     �\@      $@      �?      C@     �J@      @       @     �Q@      �?     �Q@      8@     @R@     �C@      @       @     �M@     �T@      @      $@     �P@      <@     �G@     @P@     @T@      S@      @             �H@      a@      @      &@     �V@      "@     0s@      8@      o@      O@      �?              F@      a@      �?      $@     �U@      @      s@      4@     �n@     �N@      �?              @               @      �?      @      @      �?      @      @      �?              ,@      \@     �e@      ,@      7@     �_@      0@     0q@      Q@     �h@     �\@      "@      @     �@@      J@      �?      @     �B@      @     ``@      5@     �T@     �@@              @      7@      5@      �?      @      =@      @      K@      $@      >@      ;@                       @      $@      �?              0@       @      ;@       @       @      &@              @      .@      &@              @      *@      @      ;@       @      6@      0@                      $@      ?@               @       @             @S@      &@      J@      @                      @      0@                                     �C@      @      2@      @                      @      .@               @       @              C@      @      A@      @              &@     �S@      ^@      *@      2@     @V@      &@      b@     �G@     �\@     �T@      "@       @     �P@     @W@      $@      (@      R@      $@      a@      C@     @X@     @Q@      "@      @      J@     �V@      $@      "@     �P@      $@     �Z@     �A@      W@     �M@      "@      @      .@      @              @      @              >@      @      @      $@              @      (@      ;@      @      @      1@      �?       @      "@      1@      *@                      �?      @               @      @              @      @      �?       @              @      &@      6@      @      @      $@      �?      @      @      0@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Z�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @Y3�j�C@�	           ��@       	                    @'�����@�           4�@                           �?��TXǡ@Y           ��@                          �>@���#t@           Py@������������������������       ������m@�            �w@������������������������       �°���@             :@                          �<@s�/==4	@U           ��@������������������������       �ح�� 	@           ȉ@������������������������       ��e����@;            �V@
                          �5@^7P@�           ĕ@                          �4@��@l@D           Ћ@������������������������       ��OyQ�@�           �@������������������������       �z�	�� @^            �b@                          �6@����E%@>           p@������������������������       ��K#�Fw@:            �V@������������������������       �.���]@           �y@                           @��{Pa	@�           ��@                          �3@�kR��@'           �@                           �?�9`s�@�            �q@������������������������       �!�/��@�             k@������������������������       ��R칱Q@)            �P@                           �?n��4	@s           0�@������������������������       ����`y	@7           H�@������������������������       �-��@<            @W@                           @���,�@�            �r@                           �?5.r�@_            `b@������������������������       ���לf@�?D            @Y@������������������������       ��ԓ��@             G@                           �?�ud�@_            `c@������������������������       �7�|��\@(            �O@������������������������       �՘9�9@7             W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     r@     P�@      ?@     �F@     P|@     @W@     ��@     `i@     �@      w@      <@      &@     �h@     0y@      .@      7@     0s@     @P@     @�@     �`@     (�@     �n@      4@      $@      \@      i@      @      3@     @h@     �J@     �k@     �[@     �m@     �a@      .@      �?     �F@      L@              @     �H@      @     @W@      2@     �Z@      9@      �?      �?      E@      L@              �?      G@      @     �V@      $@     �Y@      7@      �?              @                      @      @               @       @      @       @              "@     �P@      b@      @      .@      b@     �G@      `@     @W@     �`@     �\@      ,@       @     �N@      b@      @      *@     @`@      @@     �^@      T@     �^@      W@      ,@      �?      @      �?               @      .@      .@      @      *@      "@      7@              �?      U@     @i@      "@      @     @\@      (@     X�@      8@     `s@     �Z@      @             �F@      a@      @       @     �K@      @     �w@      @     @j@      G@       @              D@     �Y@      @       @     �D@      �?     �t@      @     @e@      D@      �?              @      A@                      ,@      @      G@              D@      @      �?      �?     �C@     �P@      @       @      M@      @     `b@      1@      Y@      N@      @              "@      $@      �?              (@      �?     �B@              @      *@              �?      >@      L@      @       @      G@      @     �[@      1@     @W@     �G@      @      $@     @W@     �f@      0@      6@     @b@      <@     pq@      Q@     �k@      _@       @      $@     �T@      d@      ,@      0@     @_@      ;@     �b@     �N@     `a@     @Z@       @      @      3@      B@              @      :@      @      S@      ,@     �N@     �A@              @      0@      9@               @      8@      @      I@      "@     �I@      <@                      @      &@              @       @              :@      @      $@      @              @     �O@      _@      ,@      &@     �X@      4@     �R@     �G@     �S@     �Q@       @      @      I@      [@      *@      &@     �T@      4@      L@      F@      Q@      K@       @              *@      0@      �?              0@              2@      @      $@      0@                      &@      7@       @      @      5@      �?      `@      @     �T@      3@                      @       @              @       @      �?     @S@      @     �@@      @                      @      @               @      @              O@              9@       @                       @      @              @      @      �?      .@      @       @      �?                      @      .@       @      �?      *@              J@              I@      0@                              @       @              @              1@              8@      &@                      @      "@              �?      $@             �A@              :@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�G�R@p	           ��@       	                    �?�"��@M           ��@                           �?�n7�+ 	@�           Ę@                           �?�E�z�@           �z@������������������������       ���&s@f             d@������������������������       �����@�            �p@                          �8@�ied%�	@�           �@������������������������       ���;s�@�           ��@������������������������       �[��.
@�            �v@
                           @���� �@v           h�@                           �?��5rB^@S           ��@������������������������       �r��-@�            �m@������������������������       ������`@�             s@                            �?�"{��@#             G@������������������������       �����@             0@������������������������       ��c@             >@                           �?HsU��@#           ,�@                          �4@��]�� @]           ��@                          �1@dԎ
�?�            �v@������������������������       ��g���?^            �c@������������������������       ���u���?v            �i@                          �>@�KJ��@�            �h@������������������������       ���`��r@�            `g@������������������������       ��}�F��?             &@                           @�:��d�@�           d�@                          �5@���N~n@�           �@������������������������       ���n@�           ��@������������������������       �NϞ�n�@           @|@                           7@tC�y��@             =@������������������������       ����L&@             1@������������������������       ��[���@             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      r@     (�@      <@     �L@     �{@     @T@     ��@     �g@     8�@     �u@      =@      .@     �j@     `u@      2@     �F@     @s@     �P@     �x@     �c@     �v@     �l@      6@      .@      d@     �p@      1@      B@     �m@      L@     �l@      ]@     0p@     �e@      4@              C@     �P@      �?      "@      M@      @      V@      5@     �W@     �F@      �?              ,@      1@                      3@              H@      @     �D@      1@      �?              8@     �H@      �?      "@     �C@      @      D@      1@      K@      <@              .@     �^@     �h@      0@      ;@     �f@      I@     �a@     �W@     �d@      `@      3@       @     �U@      a@      "@      5@     ``@      ;@      ]@     �H@      _@      S@      @      @      B@      O@      @      @     �H@      7@      9@      G@      D@     �J@      (@             �I@     �S@      �?      "@     �Q@      &@     �d@      E@     �Z@      K@       @              G@     �R@      �?      @     �P@      @     �c@      ?@     �X@      J@       @              2@      B@              �?      <@      @     @P@      ,@     �G@      9@      �?              <@      C@      �?      @      C@      @     �W@      1@     �I@      ;@      �?              @      @               @      @      @      @      &@       @       @                      �?      @                              @      @      @               @                      @      �?               @      @              @       @       @                      @     �S@     �i@      $@      (@     �`@      ,@     (�@      @@     �{@     �^@      @              .@      L@       @       @      9@      @      r@      "@     @a@      2@       @               @      =@               @      .@             �j@      @     �T@       @       @              �?      ,@               @      "@             �W@              A@       @       @              @      .@                      @             �]@      @     �H@      @                      @      ;@       @              $@      @     @S@      @     �K@      $@                      @      ;@       @              "@      @     �R@      @      K@      @                                                      �?              @      �?      �?      @              @     �O@     �b@       @      $@     @[@      "@     0x@      7@      s@      Z@      @      @     �M@     �b@       @      @     @Z@      @     �w@      5@     �r@      Z@      @              9@     �T@      @      @      M@      �?     �p@      *@     �h@      D@      @      @      A@     @Q@       @       @     �G@       @     �\@       @      Z@      P@       @              @                      @      @      @      @       @      @                                                      @       @      @      @              @                              @                               @      �?      @       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ3@�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @2��EE@�	           ��@       	                   �5@31[���@w           \�@                            �?4JQ6x'@�           ��@                           @�u���@�             s@������������������������       �B�P���@a            �a@������������������������       �5&Ty�@f            `d@                            �?��{ց@�           h�@������������������������       ����`�,@�            �q@������������������������       �h�%i�@=           0@
                           �?,f*�y�	@�           ��@                          �:@�S�d;	
@'           `�@������������������������       �L0'JbB	@U           @�@������������������������       �V�,>
@�            @t@                           �?f�<�@�            0p@������������������������       ��?LѴ�@(            @Q@������������������������       �A_F��@u            �g@                           @[���o�@3           l�@                           �?δ)�@�           ��@                          �4@R_����?�             w@������������������������       �3���v�?�             p@������������������������       ���~#�@J            �\@                           @oU����@           ��@������������������������       ��W��U@.           p}@������������������������       �y`��]@�            �u@                           �?��N���@A           p@                           >@REj�~�@|            �g@������������������������       �:8ND��@u            @f@������������������������       �XL��J@             *@                          �3@
�S]�@�            �s@������������������������       �u~�O�@D             \@������������������������       ���2%�@�             i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `s@     (�@      ;@      K@     0{@      U@     ��@      l@     (�@     `v@      ?@      3@     �l@     �r@      4@      D@      s@     @R@     �y@      g@     px@     `l@      ;@      @     �S@      c@      @      &@     �a@      2@     @o@     @T@     @o@      U@       @              ;@      B@              �?      ?@      @     @Q@      8@      W@      4@      @              @      ,@              �?      $@      �?      A@      @     �O@       @      �?              5@      6@                      5@       @     �A@      3@      =@      (@       @      @     �I@      ]@      @      $@      \@      .@     �f@     �L@     �c@      P@      @      @      9@     �J@       @      @      =@       @      N@      4@      I@      9@      @      @      :@     �O@      @      @     �T@      @     @^@     �B@      [@     �C@      �?      (@     �b@      b@      .@      =@      d@     �K@      d@      Z@     �a@     �a@      3@      (@     �\@     �_@      .@      6@     @`@      E@      Z@      S@     �Y@     @\@      2@              R@      W@       @      ,@     �U@      4@     �Q@      G@     �S@      I@      ,@      (@      E@     �A@      @       @      F@      6@     �@@      >@      8@     �O@      @             �B@      2@              @      ?@      *@      L@      <@      C@      >@      �?              $@       @                      @       @      <@      @      ,@      @                      ;@      0@              @      ;@      &@      <@      8@      8@      9@      �?      �?     @T@     �k@      @      ,@     ``@      &@     ��@     �C@     �{@     ``@      @      �?     �K@     �c@      �?      @     �S@      @     �}@      7@     `s@      S@       @              *@     �E@                      (@      @      h@      @      V@      ,@                      @      7@                      @             �b@      �?     �O@      @                      @      4@                      @      @     �E@       @      9@      @              �?      E@     �\@      �?      @     �P@      @     pq@      4@     �k@      O@       @      �?      B@     �N@      �?      @      J@      @      b@      .@     �[@     �E@       @              @     �J@               @      .@             �`@      @      \@      3@                      :@     �O@      @      "@      J@      @     �`@      0@      a@     �K@       @              @      :@               @      $@      �?     �Q@       @      I@      1@      �?              @      8@               @      "@             �Q@      @      H@      *@      �?                       @                      �?      �?              @       @      @                      4@     �B@      @      @      E@      @      P@       @     �U@      C@      �?              @      (@      @              0@              ?@      �?      D@      @                      1@      9@       @      @      :@      @     �@@      @      G@     �@@      �?�t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$�@ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@$�Y�!@�	           ��@       	                    �?ma�	3d@e           J�@                            �?��i���@{           8�@                          �1@��˭�@a           (�@������������������������       �"�"4�2@i             f@������������������������       �$���|�@�            Py@                           �?� ڬ$@           �|@������������������������       ��a@_             a@������������������������       ����헋@�            t@
                           �?�W�sީ@�           \�@                           �?3�i�Z�@�            �u@������������������������       �R�[@N@U            @`@������������������������       ����� @�            �j@                           @��_�@           ��@������������������������       �}��jJ@g            �d@������������������������       ���4+l�@�           Ȅ@                           �?�_���@,           ��@                           �?�B���@           �|@                            �?C�v�t@�            �j@������������������������       ��'$۝@Q            �_@������������������������       �d�0PJN@7            @U@                           @d<-!ż@�            �n@������������������������       �
�,�@/             R@������������������������       �A/"�@f            �e@                           @#�e��@           p�@                           @�KQx�l	@            �@������������������������       ��g�L	@�           ��@������������������������       �p��.�H@I            �Z@                           �?{ 2��@           �y@������������������������       �:���}@~             h@������������������������       ��ʄ�,�@�            �k@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     0t@     0�@      9@      J@     �|@      N@     ��@      j@     ��@     0w@      ?@      @      `@      s@      $@      8@     �k@      2@     (�@     @W@     �~@      d@      (@      @      J@      `@      @      *@     �]@      @     �x@      D@      i@     @R@       @      �?      9@     �W@      @      $@      R@      @     @j@      ;@      X@     �B@       @      �?      @      7@              @      .@      �?     �T@      @      ;@      (@                      5@      R@      @      @     �L@       @      `@      5@     @Q@      9@       @      @      ;@      A@      @      @      G@      @     �f@      *@      Z@      B@              @      1@      *@       @      �?      <@      @      ?@      @      6@      (@                      $@      5@      �?       @      2@      �?      c@      $@     �T@      8@               @     @S@      f@      @      &@     @Z@      &@     �u@     �J@     r@      V@      $@              0@     �J@              �?      :@              `@      "@     @W@      0@       @              &@      >@              �?      .@              =@      @      ;@      &@                      @      7@                      &@             �X@      @     �P@      @       @       @     �N@      _@      @      $@     �S@      &@     �k@      F@     �h@      R@       @       @      4@      2@              @      8@      @     �@@      *@      A@      &@      @             �D@     �Z@      @      @     �K@      @     `g@      ?@     @d@     �N@      @      "@     @h@     @q@      .@      <@      m@      E@     �q@      ]@     Pq@     @j@      3@      �?     �C@      U@               @      I@       @     �Y@      .@     @W@     �I@      @      �?      ?@     �F@               @     �A@      �?      ;@       @      @@      6@       @      �?      1@      :@              @      0@      �?      4@      @      7@      *@       @              ,@      3@              @      3@              @      @      "@      "@                       @     �C@                      .@      @     �R@      @     �N@      =@      @              @       @                      @      �?      8@      @      .@      @      @              @      ?@                      &@      @     �I@      �?      G@      6@               @     `c@      h@      .@      4@     �f@      A@     `f@     @Y@      g@     �c@      ,@       @      ^@      `@      .@      .@     @_@      >@     �Q@     �T@      X@      `@      *@      @     �Y@      [@      *@      .@     @[@      ;@      Q@     �N@     �V@     �]@      $@      @      2@      5@       @              0@      @      @      5@      @      $@      @             �A@     �O@              @      M@      @      [@      3@      V@      ?@      �?              .@     �D@              @      0@       @      J@      @     �E@      (@      �?              4@      6@              �?      E@       @      L@      *@     �F@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJi�`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��K�OJ@�	           ��@       	                    @V�6��@Y           �@                           �?"����@�           ��@                           @�8�"@�           ��@������������������������       �c���K@�            @u@������������������������       �A`Y��T@�            @x@                          �3@0^8@�            �t@������������������������       ��*Q�j@�            �i@������������������������       ���q��@R            �^@
                           @��l�̾@�           ��@                           @�o��\@�            �q@������������������������       ��<�>�@�             m@������������������������       �����W@             I@                            �?��so�@           0�@������������������������       �:�8��^�?s            �h@������������������������       �ܑq��@�           �@                           �?v���ө@M           �@                          �<@I�u6�@&           p~@                           �?`�H[� @�            �v@������������������������       ����a@f            `c@������������������������       �G��߿h@�             j@                           @;�C�4�@>             _@������������������������       �0���%@,            @T@������������������������       �'ޤ�7 @            �E@                          �=@���0	@'           ��@                          �7@b%{�	@�           ܐ@������������������������       ���T�@           �w@������������������������       ��R�-7*	@�           Ѕ@                           �?Y���y�@h             e@������������������������       �A\��%@!             J@������������������������       ��Lb(Ō@G            @]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@      �@      ;@     �O@     �{@     �R@     ��@      k@     ��@     `w@      =@      @     �`@     r@      *@      @@     �l@      5@     ��@      W@     �}@      f@      &@      @     @T@     �c@      $@      4@     `b@      ,@     `l@     �S@     �h@     �\@       @      @     @Q@     �X@      @      ,@     �Y@       @     �`@     �M@      a@      W@       @      @      ?@      C@       @      @      B@       @      T@      >@     @S@      A@      @              C@     �N@      @      $@     �P@      @      J@      =@      N@      M@      @              (@      M@      @      @     �F@      @     �W@      3@     �N@      6@                      $@      @@              @      6@      @     �P@      (@     �D@      1@                       @      :@      @      @      7@      @      =@      @      4@      @                     �J@     �`@      @      (@     @T@      @     �}@      ,@     `q@     �O@      @              :@      C@                      6@      @     @Y@      @      O@      5@      �?              2@      @@                      6@      @     �T@      �?     �L@      0@                       @      @                              �?      3@      @      @      @      �?              ;@     �W@      @      (@     �M@      �?     `w@       @      k@      E@       @               @      0@              �?      7@              Z@             �G@      @                      9@     �S@      @      &@      B@      �?     �p@       @      e@     �C@       @      *@     �f@     �o@      ,@      ?@     `k@      K@      t@     @_@     @s@     �h@      2@       @      C@     @S@      @      @     �L@      @     @_@      ;@     @Y@     �D@      @       @      ?@     �P@      @      �?     �E@      @     @X@      1@     �S@      1@      �?       @      9@      >@       @      �?      <@       @      5@      "@      <@      @      �?              @     �B@       @              .@       @      S@       @     �I@      &@                      @      $@              @      ,@       @      <@      $@      6@      8@       @              @      @              @      *@               @      "@      $@      7@       @                      @                      �?       @      4@      �?      (@      �?              &@     �a@     @f@      $@      9@     @d@      H@     `h@     �X@     �i@     �c@      .@       @      ^@     �b@      $@      9@     �a@     �D@      f@     �T@      h@     �]@      ,@      @     �J@      Q@      @      $@      E@      &@      R@      5@      M@      B@      @      @     �P@     �T@      @      .@      Y@      >@      Z@     �N@     �`@     �T@      &@      @      7@      <@                      4@      @      3@      0@      ,@      C@      �?      @       @      $@                      $@      @      @      @      @      @                      .@      2@                      $@      @      *@      *@      $@      A@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJHž\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�@q|�@�	           ��@       	                   �2@��F�@v           L�@                           �?��V�v@�           X�@                           �?n���'@(           �~@������������������������       ��6 �7D@�            @m@������������������������       ����0��@�             p@                           �?�}@��t@`           `�@������������������������       �Ft�R<@�             j@������������������������       ���@f��@�            �u@
                            �?�&x@��@�           �@                            �?���e�@           z@������������������������       ��)����@~             h@������������������������       ����@�             l@                           @�"��@�            �u@������������������������       �L���N@�             m@������������������������       ��&�駙@L             ]@                          �;@�d}���@<           l�@                           @R��*7@           x�@                           �?�^�14	@l           ��@������������������������       �_���^	@�            `u@������������������������       �EQB��@�           0�@                           @T"�D�@�           �@������������������������       �J�g���@�           ��@������������������������       �mwc���@)            �P@                           �?�O"���@!           �}@                           �?',���@�            `q@������������������������       �Y�fʉ�@>            �Y@������������������������       ��D��;	@m            �e@                           @�MbrT@v            @h@������������������������       ���ҿ�B@3            �U@������������������������       �,�O�@�@C            �Z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     0s@     @�@      :@     �L@     �y@     �W@     ؎@      n@     ��@     `x@      @@      @     @Y@     Pp@      @      3@      c@      0@     P�@     �V@      w@     @d@      (@      �?      M@      d@      �?      @     @V@      @     py@      F@      g@     �T@      @      �?      8@     �S@      �?      @      J@      @     `h@      .@     @R@     �E@                      $@      <@              �?      8@      �?     �^@       @      >@      0@              �?      ,@     �I@      �?       @      <@      @     @R@      *@     �E@      ;@                      A@     @T@              @     �B@       @     �j@      =@     �[@     �C@      @              &@      7@                      $@              [@      @     �C@      $@      @              7@      M@              @      ;@       @      Z@      8@      R@      =@      @      @     �E@     @Y@      @      (@     �O@      $@     `j@     �G@      g@      T@      @              ;@      F@      @       @     �C@      �?     �Z@      =@     @\@      H@       @              &@      0@                      5@              J@      3@     �L@      .@       @              0@      <@      @       @      2@      �?     �K@      $@      L@     �@@              @      0@     �L@      �?      $@      8@      "@      Z@      2@     �Q@      @@      @       @      .@      F@              @      0@       @     @S@      @     �E@      6@      �?      �?      �?      *@      �?      @       @      @      ;@      .@      <@      $@       @      1@     �i@     0r@      3@      C@      p@     �S@     w@     �b@     �z@     �l@      4@      @     `c@     @m@      .@      =@     �h@     �L@     0t@      [@     pv@      `@      3@      @     @_@     �a@      "@      6@     �`@     �@@     �_@     �U@     `f@     �S@      .@      �?     �E@      H@      @      "@      D@      &@     �L@     �@@     �K@      @@      "@      @     �T@      W@      @      *@     �W@      6@     �Q@     �J@      _@     �G@      @      �?      >@     �W@      @      @     �N@      8@     �h@      6@     �f@     �H@      @      �?      8@      U@      @      @      L@      4@      g@      &@     @e@     �G@                      @      $@      @              @      @      (@      &@      $@       @      @      $@     �I@     �L@      @      "@      O@      6@      G@     �D@     @Q@      Y@      �?      $@      ?@     �@@      @      @      @@      3@      ,@      9@      ;@     �S@      �?      @      "@      3@              �?      .@       @      @      @      "@      ?@              @      6@      ,@      @      @      1@      &@      &@      4@      2@     �G@      �?              4@      8@              @      >@      @      @@      0@      E@      6@                      @      .@              @      @       @      2@      .@      ,@       @                      1@      "@                      7@      �?      ,@      �?      <@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ.�(WhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @>>�~h@�	           ��@       	                    �?��0��@�           ȡ@                          �6@�:U]�@�           ��@                            �?da$ooV@�            Pz@������������������������       ���Eۃ�@I            �_@������������������������       ��{9?�@�            pr@                           �?�	m�Nc@�            �p@������������������������       ��
�@�             k@������������������������       ��4���@            �I@
                           �?4��SN	@�           ̘@                          �4@��ny�	@�           �@������������������������       ��2}k�@           �{@������������������������       �U���z�	@�            �@                            �?�z+|��@
           �{@������������������������       ��{��;�@M             a@������������������������       �h�K;z@�             s@                          �3@0A��J@            ��@                           �?�t|�Ѡ@�           ��@                          �2@a\�| ��?�            0r@������������������������       �x�_���?�            @l@������������������������       ��V�Y�?#            @P@                            �?���ó�@           �y@������������������������       ����c@>            �V@������������������������       �ɖ�9�@�             t@                          �=@�e���@N           8�@                           @PݘKM@*           p�@������������������������       ������P@f           ��@������������������������       ���g���@�            �s@                           @��s�TJ@$            �L@������������������������       �ޯ5��@             ;@������������������������       �!`��x@             >@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@      r@      @      A@      O@     ~@     @T@     <�@      l@     �@     �u@      >@      9@     �j@     Pt@      9@      G@     �t@     �J@     �y@     `f@     �x@     �m@      :@      @     �P@     @U@      @       @     @U@       @     @e@      B@     �c@      L@      @              E@     �G@              @      D@      @     �_@      4@     �[@      7@      �?              $@      .@              �?      @      @      C@      �?     �G@      @                      @@      @@              @     �@@      @      V@      3@     �O@      4@      �?      @      9@      C@      @      @     �F@      �?      F@      0@     �H@     �@@      @      @      8@      @@      @      @      D@      �?      8@      .@      B@      ?@      @              �?      @                      @              4@      �?      *@       @      @      5@     �b@      n@      5@      C@      o@     �F@     �n@     �a@     �m@     �f@      3@      5@     �\@     �c@      3@      7@     `h@     �B@      b@     @[@     �d@      b@      2@      @      @@     �D@      @      @     �S@      *@      S@     �@@     @T@     �O@      @      .@     �T@     �]@      (@      0@     @]@      8@      Q@      S@     �T@     @T@      (@              A@     @T@       @      .@     �J@       @     @Y@      A@      R@     �C@      �?              @      2@              @      *@      @     �E@      $@      5@      0@      �?              <@     �O@       @      &@      D@      @      M@      8@     �I@      7@              @     @R@     �e@      "@      0@     �b@      <@     ��@     �F@      y@      \@      @              =@     �Q@      @      @      C@      �?      u@      ,@      e@      B@      �?              @      7@                      $@             �e@      @     �P@      $@      �?              @      1@                      @             `a@      @      G@      $@      �?                      @                      @             �A@              4@                              9@     �G@      @      @      <@      �?     @d@      &@     �Y@      :@                       @      *@                      @              F@      @      ,@      &@                      7@      A@      @      @      8@      �?     �]@       @      V@      .@              @      F@     �Y@      @      $@     �[@      ;@      r@      ?@     @m@      S@      @      @      C@     �W@      @       @     @X@      :@     �q@      :@     `l@     �P@      @      @      =@     �K@              @     �M@      (@     �h@      &@      c@     �D@       @              "@      D@      @      @      C@      ,@     �U@      .@     �R@      :@      �?              @       @       @       @      *@      �?      @      @      @      "@                      @      �?               @      @              �?      @      @      @                       @      @       @              "@      �?      @       @       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��IhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                              @� �Q>B@�	           ��@       	                    �?s#Zj�@�           ڥ@                           �?j����@=           8�@                            �?�d��@           �{@������������������������       �M�u���@b             c@������������������������       ��S]�l:@�            Pr@                          �4@�8�Gx�@#           �|@������������������������       ��u�P �@�             p@������������������������       ��`x>��@�            �h@
                           @MT$�@�           ��@                          �4@u\2S�/	@8           (�@������������������������       �F�,g��@�            Pv@������������������������       ����k	@V            �@                           �?͊��X@l           �@������������������������       �m���@-           `~@������������������������       �V��|@?           �@                          �3@N{�2:@�           p�@                           �?��uԝ�@�            �v@                          �0@G?5��A@s             h@������������������������       �ʿ��i��?             .@������������������������       �$�v�,h@k             f@                           @;9��
@h             e@������������������������       �
�Ӳ�?1             T@������������������������       �ד�u�@7            @V@                          @@@Q|Pn��@�           ��@                           @z!��ժ@�           ��@������������������������       ��^�c �@r           ��@������������������������       ������@O            �`@������������������������       �'tdX@             >@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     `r@     0�@      @@     �M@     {@     �U@     ��@     `k@     �@     0u@      @@       @     �i@     �w@      *@      E@     �q@      N@     ȇ@      c@     ��@     �m@      2@      �?      N@      `@       @      @     @S@      @      t@      :@     @l@     �H@      @      �?      :@     �L@               @      @@      @     `f@      0@     �W@     �@@      �?      �?      �?      1@                      2@       @     @Q@       @      @@      &@                      9@      D@               @      ,@       @     �[@      ,@     �O@      6@      �?              A@      R@       @      @     �F@      �?     �a@      $@     ``@      0@       @              5@      H@                      *@              Z@      @     �I@      *@      �?              *@      8@       @      @      @@      �?     �B@      @      T@      @      �?      @      b@     �o@      &@     �B@     @j@     �K@     �{@     �_@     Py@     �g@      .@      @     �T@     �`@      @      2@     �`@     �E@     @^@     �X@     �a@      [@      *@      �?      8@     �E@      �?      @     �N@      @     �R@     �C@      M@      D@       @      @     �M@     @V@      @      *@     @R@      D@     �G@      N@     �T@      Q@      @      �?     �N@     �^@      @      3@      S@      (@      t@      <@     �p@      T@       @      �?      8@      P@       @      ,@      F@      @      c@      ,@     �]@      F@       @             �B@      M@      @      @      @@      @     �d@      ,@     @b@      B@              &@     �V@     �`@      3@      1@     @b@      ;@     �o@     �P@     �m@     �Y@      ,@      @      7@      D@       @      @      E@       @     �_@      (@     �R@      4@              @      *@      6@       @      @      A@       @     �E@      @      B@      .@                              �?                      &@              �?      �?      �?                      @      *@      5@       @      @      7@       @      E@      @     �A@      .@                      $@      2@              �?       @             �T@      @     �C@      @                      �?      @              �?                     �I@      @      .@      @                      "@      .@                       @              @@      �?      8@                      @     �P@     �W@      1@      &@      Z@      3@     �_@      K@      d@     �T@      ,@      �?     �P@      W@      1@      &@     @X@      3@     �_@      I@     �c@     �R@      ,@      �?     �O@     @V@      *@      @     @V@      0@      T@     �F@     @^@      L@      ,@              @      @      @      @       @      @      G@      @     �A@      3@              @              @                      @              �?      @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?߉��A@�	           ��@       	                    �?���/@           h�@                          �7@��3@�           ��@                           @��x�@2           P~@������������������������       �y#�K@@�            �p@������������������������       ���H��?�             k@                          �>@����t@h            �e@������������������������       ����!B@[            �b@������������������������       �pC�#$@             6@
                            �?+��Ŧ�@x           H�@                          �4@��l��@�            �t@������������������������       ����V��?k            `d@������������������������       ��
0_@f             e@                          �1@�D��P�@�            �o@������������������������       �Ը��k��?'            �P@������������������������       ���x��@�            `g@                           �?)�(�=E@�           ޤ@                           @`Y��U	@x            @h@                           �?�)�Md	@_            `c@������������������������       ���Ɏ�@7             V@������������������������       �!��X/	@(            �P@                            �?�����@            �C@������������������������       �y���@             9@������������������������       ���h%vO@             ,@                           @8�/��@>           Z�@                          �5@&�e�&�@u           �@������������������������       ���D��M@�           p�@������������������������       ���4G�@�           (�@                           �?8��R+	@�            �r@������������������������       �-ޙ��5	@Q            �]@������������������������       ���.P�@x            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     r@     ��@      ;@      P@     `|@     @T@     H�@     �k@     �@      v@      ?@      �?     @R@     �e@      @      ,@     �Z@       @     �}@      D@     0q@      Q@      @      �?     �@@     �V@      @      &@      M@      @     �p@      3@     �_@      C@      �?              0@     �Q@      �?      @      G@      @     �j@      ,@     @W@      3@      �?              ,@      H@      �?      �?     �A@      @     �U@      ,@      I@      *@      �?               @      7@              @      &@             �_@             �E@      @              �?      1@      4@       @      @      (@       @      K@      @      A@      3@              �?      (@      4@       @      @      &@             �H@      �?      @@      1@                      @                      �?      �?       @      @      @       @       @                      D@      U@              @      H@      �?      j@      5@     �b@      >@       @              5@      J@                      4@              \@       @      Z@      (@       @               @      6@                      @             �R@              I@      @                      *@      >@                      .@              C@       @      K@       @       @              3@      @@              @      <@      �?      X@      *@      F@      2@                      @      @                      @              D@       @      (@                              0@      <@              @      6@      �?      L@      &@      @@      2@              ,@      k@     px@      8@      I@     �u@     @R@     ��@     �f@     �~@     �q@      <@      @      .@      6@              "@     �A@      @      1@      ;@     �B@      1@      @      @      &@      6@              "@      @@      @      $@      4@      :@      &@      @       @       @      $@               @      4@      �?      @      &@      4@      @      @       @      @      (@              @      (@      @      @      "@      @      @                      @                              @      �?      @      @      &@      @                                                      @              @      @       @      @                      @                                      �?      �?      @      @       @              $@      i@     w@      8@     �D@     �s@     �P@     (�@      c@     �|@     �p@      7@      @     �d@     �t@      8@      C@     0q@      H@     �~@     @^@     Pz@      n@      0@      @      O@     �h@      @      ,@     �]@      .@     @t@      O@     p@     @\@      @      @     �Y@     �`@      1@      8@     �c@     �@@     �d@     �M@     �d@     �_@      $@      @      B@     �B@              @      C@      3@      M@      @@     �B@      =@      @      @      .@      *@                      4@      (@      3@      1@      @       @      @              5@      8@              @      2@      @     �C@      .@      ?@      5@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ɃhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�^�9@�	           ��@       	                   �;@Vz��n4	@�           �@                           @�����@J           ��@                           �?�eE��~@9           ��@������������������������       ��9`I@2           �~@������������������������       ��3���@           ��@                          �5@%̓P2@             =@������������������������       ��g�L@             *@������������������������       �����@	             0@
                          @@@�U��4�	@�             p@                           @��u��2	@�             k@������������������������       �ѕr�M�@^            `c@������������������������       �סMXP@$             O@                          �@@g_&>��@            �D@������������������������       �|R��>@	             0@������������������������       ������@             9@                            �?�ω`�@�           �@                           @F[����@1           ��@                           @�)YɁ@�           D�@������������������������       ��+a~�@D            ~@������������������������       ��s��@�           x�@                          �6@J�\�@<            �U@������������������������       �����@%             L@������������������������       �I��@             >@                           �?1k8H�@�           ��@                          �3@�9��@-           @~@������������������������       ��4N:� @�            �i@������������������������       ��)כ�@�            Pq@                           @�n�+��@c           �@������������������������       �Q�i��@           �{@������������������������       �3�k9�@R            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �s@      �@      8@      H@     P|@      W@     ��@     �l@     8�@     �u@      =@      *@     �i@      m@      1@     �@@     �m@     �J@     @k@      b@     �p@      d@      7@      "@      f@      h@      (@      ;@     �h@      =@     @i@     @_@      n@     �\@      3@      @     �e@     �g@      (@      ;@     `h@      <@      i@     �^@      n@     �[@      $@             �G@     @Q@      �?      (@     �T@      "@     �Z@      ?@      W@      F@      �?      @     @_@     @^@      &@      .@     @\@      3@     �W@     �V@     �b@     �P@      "@      @      @       @                       @      �?       @      @              @      "@      @       @                                      �?       @                       @      @               @       @                       @                      @              �?      @      @      <@      D@      @      @      E@      8@      0@      3@      7@     �G@      @       @      :@      >@      �?      @      A@      7@      0@      1@      1@     �E@      @       @      8@      >@      �?      @      7@      &@      (@       @       @      >@      @               @                      �?      &@      (@      @      "@      "@      *@      �?       @       @      $@      @       @       @      �?               @      @      @                       @       @      @              �?                              @      �?               @               @               @      @      �?               @              @                     �[@     �s@      @      .@     �j@     �C@     ��@     @U@     ��@     �g@      @             �R@      e@      @      "@     �Z@      5@     �y@      F@     ps@      Y@      �?             �P@     �c@      @      "@     �Y@      0@     �x@      A@     �r@      U@      �?              <@     @R@      �?      @     �I@      &@     @a@      3@     @]@     �C@      �?             �C@     �T@      @      @      J@      @     �o@      .@     @g@     �F@                      @      *@      �?              @      @      7@      $@       @      0@                      �?      $@      �?              �?      @      6@      @      @      &@                      @      @                       @      �?      �?      @      @      @                     �B@     �a@       @      @      [@      2@     �w@     �D@      m@      V@      @              $@     �M@       @       @      E@      @     �g@      6@     @Y@      I@      �?              @      9@                      *@              Z@      "@     �E@       @                      @      A@       @       @      =@      @      U@      *@      M@      E@      �?              ;@      U@              @     �P@      &@     �g@      3@     ``@      C@      @              3@     �O@              @      D@      $@     �c@      .@     �W@      B@      @               @      5@                      :@      �?      ?@      @      B@       @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���7@�	           ��@       	                    �?VG}#@�           0�@                          �1@0�ʡ@�           �@                          �0@��27	- @�             r@������������������������       ���ܠ� @A             Y@������������������������       ���4P���?u            �g@                           �?��Vg�@�            �w@������������������������       ���A(�y@Y            �`@������������������������       ��=6�;@�             o@
                           @���g�L@�           ��@                          �3@�%��@�           ��@������������������������       �M\X@O           @�@������������������������       ����(�@u            �f@                          �3@Q��' ^@"           �|@������������������������       ���'��/@�            0v@������������������������       ��Kq�T�@B             [@                           @CJ��5�@           ��@                           �?� ��Af	@5           d�@                          �;@^��*o@�            @v@������������������������       ��P:��@�            �p@������������������������       ���Bћ%@8            �V@                            @�dA��	@K           ��@������������������������       �yC<Sj	@c           ��@������������������������       ������	@�            �w@                           @@҄�Wq@�            �@                           @�ʣY�@M           �@������������������������       ��N`�ɵ@�            �t@������������������������       ��&�#N*@z            �e@                           @�����k@�            �l@������������������������       ��9/u�@�            `j@������������������������       ���֣�@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pr@     ��@      B@      C@     �|@     @X@     ��@     �i@     0�@     �t@      <@      @     �X@     �o@       @      2@      f@      :@     ��@     @U@     0{@      ^@      @              =@     �S@              @      F@      @      r@      5@     �d@      C@      �?              "@      :@                      8@             �b@      @     @Q@      "@      �?                      (@                      &@             �H@       @      6@      @                      "@      ,@                      *@             �X@       @     �G@      @      �?              4@     �J@              @      4@      @     �a@      1@     �X@      =@                      "@      9@                      (@      @     �@@      @      @@      .@                      &@      <@              @       @             �Z@      &@     �P@      ,@              @     �Q@     �e@       @      .@     �`@      7@     �u@      P@     �p@     �T@      @      @     �K@      [@      @      "@     �Y@      6@     `e@     �L@     ``@      O@      @      @      F@     @S@      �?      @     �M@      0@     `b@     �F@      Y@      I@      �?              &@      ?@      @       @      F@      @      8@      (@      ?@      (@      @              .@     �P@      @      @      =@      �?     `f@      @      a@      4@                      (@     �D@      @      @      <@              a@      @     �[@      0@                      @      9@               @      �?      �?      E@      @      ;@      @              1@     �h@     �s@      <@      4@     �q@     �Q@      x@     �]@     0w@     �j@      7@      .@      d@     �i@      9@      1@     �i@      K@      d@     �X@     �g@     @c@      2@      �?      D@     �L@      @      @     �J@      @     �R@      .@     �Q@      <@      @              @@      B@      @      �?      D@      �?     @Q@      "@      N@      &@      @      �?       @      5@              @      *@       @      @      @      &@      1@      �?      ,@     @^@     �b@      5@      &@      c@     �I@     �U@     �T@      ^@     �_@      ,@      @     �Q@     �S@       @       @     �W@      A@      D@     �O@     @S@      T@      @       @      I@     �Q@      *@      @      M@      1@      G@      4@     �E@      G@      @       @     �A@     @\@      @      @     �S@      1@      l@      5@     �f@     �M@      @       @      &@     �T@      �?       @      G@      *@     @f@      $@      `@     �A@               @      @     �F@              �?      ?@      $@     �`@      @     @U@      2@                      @      C@      �?      �?      .@      @      F@      @     �E@      1@                      8@      >@       @      �?      @@      @      G@      &@      J@      8@      @              6@      =@      �?      �?      9@             �E@      $@     �I@      8@      @               @      �?      �?              @      @      @      �?      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ
�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@z����s@�	           ��@       	                    @��R�*@o           $�@                            @��؎@"           H�@                           @&�R��@U           ��@������������������������       �v�	�@�             w@������������������������       ���C�K@m             d@                           �?A��L��@�            `s@������������������������       ���@8            �V@������������������������       ��]CsQ	@�            �k@
                           �?{_����@M            �@                            �?󾎧L�?�             w@������������������������       �&�SK�� @{            �f@������������������������       �\�'���?l            `g@                          �1@��˖�&@f           p�@������������������������       �K�/��< @t            @i@������������������������       ��k<"U@�            @x@                            @PD��@3           ��@                           @㶢� �@�           �@                          �:@x�¡�	@	           ��@������������������������       ��ޞJb	@h           ��@������������������������       ���� ��	@�            �o@                           @��W�t�@�           0�@������������������������       �I"��R@           |@������������������������       ��X��@�            �h@                           �?�0-�X|@�           8�@                          �8@�'�K�@b            �d@������������������������       ����E�3@5            @W@������������������������       � c�v4]@-            @R@                           �?��"Y��@4           ~@������������������������       ��K�\R�@            �E@������������������������       ��>^h�@           `{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �t@     �~@      8@      L@     �}@     �T@     ��@     �l@     `�@     �v@     �B@      @     @Z@      h@      $@      .@     `f@      2@     ��@     �S@     @z@     @a@       @      @     �N@     @W@      @      "@     @_@      .@     �h@     �M@     `e@     @V@       @      �?      <@      H@       @      @     @S@      "@     �_@     �B@     ``@     @P@      @              5@      A@              @      N@      @      U@      ,@      Z@     �E@       @      �?      @      ,@       @              1@      @      E@      7@      ;@      6@       @      @     �@@     �F@      @      @      H@      @     @R@      6@      D@      8@      @              *@      &@                      4@              6@      �?      ,@      "@              @      4@      A@      @      @      <@      @     �I@      5@      :@      .@      @              F@     �X@      @      @      K@      @      {@      3@      o@     �H@                      *@      C@              �?      *@             �j@      @     @Q@      ,@                      $@      7@              �?      $@              X@       @      ?@      $@                      @      .@                      @             �]@      @      C@      @                      ?@     �N@      @      @     �D@      @      k@      (@     �f@     �A@                       @      .@              �?       @             @V@       @      Q@      &@                      7@      G@      @      @     �@@      @      `@      $@      \@      8@              ,@     @l@     �r@      ,@     �D@     �r@      P@     �v@      c@     �x@      l@      =@       @      c@     �i@      "@      @@      h@      H@      p@     �Y@      r@     �a@      :@       @     �Y@     �\@      @      ;@     �_@     �D@     �T@     @S@     @^@     �V@      5@      �?     �S@     �V@      @      6@     �U@      6@     �Q@      K@     @U@      C@      0@      @      9@      8@      @      @      D@      3@      (@      7@      B@     �J@      @              I@     �V@       @      @     �P@      @     �e@      9@      e@      J@      @              ?@     @Q@       @      @      F@      @     �`@      3@     �[@      =@                      3@      5@              �?      7@              D@      @     �M@      7@      @      @     @R@     @W@      @      "@     �Y@      0@      Z@     �I@     �Y@     �T@      @              (@      6@              @     �A@             �E@      &@      >@      $@                      @      ,@                      (@              <@      @      6@       @                      @       @              @      7@              .@       @       @       @              @     �N@     �Q@      @      @      Q@      0@     �N@      D@      R@      R@      @       @      &@      $@                      @      @              @       @      @      �?      @      I@     �N@      @      @     �O@      *@     �N@      A@     �Q@     @Q@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�߀UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���/��@�	           ��@       	                   �1@Xm�	@|           ��@                           �?&���=@�            �r@                          �0@�Wl��L@�            �i@������������������������       �ҋ�@'             O@������������������������       ��'�er�@Z            �a@                           �?�ʃ�V� @9            �W@������������������������       �GM[A�	�?             :@������������������������       �F%��� @'            @Q@
                           �?���n7X	@�           H�@                           �?t80��	@           ��@������������������������       �A�M��(@�            �x@������������������������       �P� �
@�            �@                           �?�-�=SS@C           0~@������������������������       �n\����@a            @a@������������������������       ���ל�@�            �u@                           @*@�4@N           0�@                           �?�Fr�]@�           �@                           @~A݊�x @�            Px@������������������������       ����d5@�            Pp@������������������������       ��Ǯ S��?L             `@                          �2@-�?@           ��@������������������������       �Y#���2@�            �m@������������������������       �z��[��@f           @�@                            @M:D��@V           ��@                          �;@c���@           `y@������������������������       ��I���b@�            �v@������������������������       �+�E@            �C@                           @[B	
D�@N            �^@������������������������       �,���S1�?+            �O@������������������������       ��R8H`@#             N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@      A@     �M@     �|@     �T@     ��@      k@     ��@      x@      >@      2@     �k@     �s@      8@     �G@     s@     �P@     pu@     @f@     �v@     pp@      ;@       @      4@     �J@      �?      @      <@       @      Z@      ,@     �I@      5@               @      1@     �B@      �?      @      :@       @      M@      @      A@      2@                      @      &@              @      (@              0@       @      @      @               @      $@      :@      �?              ,@       @      E@      @      =@      (@                      @      0@                       @              G@       @      1@      @                      �?      @                      �?              (@               @      �?                       @      *@                      �?              A@       @      "@       @              0@      i@     `p@      7@      F@     Pq@      P@     �m@     �d@     �s@     @n@      ;@      0@      d@      h@      6@     �C@     `j@     �H@     `c@     @^@     @j@     �g@      ;@       @      I@      L@      @      @      C@      @     �P@      ?@      U@      H@      @      ,@     �[@      a@      3@     �@@     �e@      E@     @V@     �V@     �_@     �a@      7@              D@     �Q@      �?      @     �P@      .@      U@     �E@     �Z@     �J@                      &@      2@              �?      ,@       @     �C@      @     �D@      @                      =@      J@      �?      @      J@      *@     �F@      C@     @P@      G@                     �W@     @o@      $@      (@     `c@      0@     @�@      C@     �z@     @^@      @             �P@      f@      �?      @     @[@      &@     0|@      4@     �r@      R@      �?              ,@      E@                      =@      @     `i@      @     @T@      "@                      @      =@                      4@      @      `@      @      M@       @                      @      *@                      "@             �R@              7@      �?                      J@     �`@      �?      @      T@      @      o@      .@     `k@     �O@      �?              (@     �C@                       @      �?     �S@      �?      R@      :@                      D@     �W@      �?      @      R@      @      e@      ,@     `b@     �B@      �?              <@     �R@      "@       @      G@      @     �d@      2@     @_@     �H@       @              8@      P@      @      @     �A@      @     �\@      0@      Y@     �@@       @              2@     �K@      @      @      <@      @     �\@      ,@     �W@      ;@       @              @      "@      @              @              �?       @      @      @                      @      $@       @      @      &@              I@       @      9@      0@                       @                      @      @              B@       @      ,@      @                       @      $@       @               @              ,@              &@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ƈEhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @��
l��@�	           ��@       	                   �5@�E�u	@�           t�@                           �?��q���@�           �@                            �?��xT�@�            �w@������������������������       �DfR��@D             Z@������������������������       �Y���@�            @q@                            �?TtC��[@�            �@������������������������       �A�-W��@�            @w@������������������������       ��+��qd@�            �t@
                          �7@u !���	@�           ��@                           @��|�@�            �u@������������������������       ����y@�             i@������������������������       �ya�_�@a            @b@                          �<@<�p
@�           �@������������������������       ��w�(_{	@I           ��@������������������������       �A���%
@�            0q@                          �7@LӢs�@           <�@                           @�p��@            �@                            �?B7�<��@           ��@������������������������       �2�zh2�@�            0r@������������������������       �a��,@Z           `�@������������������������       ���x�@             1@                           �?�v�@�            �x@                           @{Ǐ��@y            �h@������������������������       �Ĩ6��@H            �]@������������������������       ��_S�e0@1             T@                           @���I��@�             i@������������������������       �{Ӟ'�@O             _@������������������������       �ng��@4            @S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     `t@     ��@      <@     �I@      {@     @V@     �@     `k@     ��@     �x@     �E@      0@     �m@      s@      3@     �D@     �s@     @Q@     0w@     `g@     `v@     �q@     �A@      @     �R@     @c@      @      (@     `b@      9@     @n@     �R@     @i@     ``@      $@              >@     �H@       @       @     �D@      @     �[@      1@     @W@      =@      �?              @      1@              �?      @             �@@      �?     �B@      @                      :@      @@       @      �?     �A@      @     @S@      0@      L@      8@      �?      @     �F@     @Z@      @      $@     �Z@      3@     �`@      M@     @[@     �Y@      "@      �?      ?@     �N@      �?       @     �I@      ,@     �R@      9@     �N@      G@      @      @      ,@      F@       @       @     �K@      @      M@     �@@      H@      L@      @      $@     @d@      c@      ,@      =@     �d@      F@      `@      \@     �c@     �b@      9@      �?      R@     �L@       @       @      H@      @      B@      6@      Q@      6@      @             �G@      :@       @      @      ;@      �?      =@       @     �G@      &@              �?      9@      ?@              @      5@      @      @      ,@      5@      &@      @      "@     �V@     �W@      (@      5@     �]@     �C@     @W@     �V@      V@      `@      3@      @     �I@     �O@      @      @     @V@      5@     �S@      K@     �O@      S@      *@      @     �C@      @@      @      ,@      =@      2@      ,@      B@      9@     �J@      @      �?     @V@     `l@      "@      $@     @^@      4@     P�@      @@      {@     �[@       @             �N@     �f@       @       @     �S@      .@     8�@      ,@     pt@     �M@       @             �N@     �f@      @       @      S@      &@     0�@      ,@      t@     �K@       @              (@     �D@      �?              6@      @     �a@       @     �J@      0@                     �H@     �a@      @       @      K@       @     �w@      (@     �p@     �C@       @                              �?               @      @      �?              @      @              �?      <@      F@      �?       @     �E@      @     �X@      2@     �Z@     �I@              �?      1@      <@              �?      ,@             �L@      @     �H@      9@              �?      @      6@              �?      @              G@      �?      ;@      "@                      &@      @                      "@              &@      @      6@      0@                      &@      0@      �?      �?      =@      @      E@      (@      M@      :@                      @      (@              �?      2@      @     �A@      @      <@      ,@                      @      @      �?              &@       @      @      @      >@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ|��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?/���"@�	           ��@       	                    �?TL�Yv@�           ؒ@                           �?�PH&@6           �~@                            �?n�`*-�@�            �l@������������������������       �p2�*:$@)            �L@������������������������       �ٿO��K@g            `e@                           �?�;e!�@�            �p@������������������������       �$v5���@F            @[@������������������������       �2��'�@`            �c@
                            �?y�g^"�@�           8�@                           @�,��2
 @v             e@������������������������       �c�7��> @J             \@������������������������       �%�X��?,             L@                          �1@��c��@S           ��@������������������������       �NbC͑�?T             `@������������������������       �JyEn5c@�            �y@                          �4@ *�XT @�           &�@                           @�w�M@�           �@                           @'�a�ȉ@�            �k@������������������������       ���h�{3@Q            @^@������������������������       �u��8T�@?            �Y@                           @dZ=�A�@P           �@������������������������       �V�&BUZ@b           0�@������������������������       �ik����@�            �w@                           �?G�B-|�@�           H�@                           @�|���@}           ��@������������������������       �[�~���	@�            `s@������������������������       �%�;�7�@�            �r@                           @��|ɞ@<           ��@������������������������       �u�A�	@�           ؃@������������������������       ��`��q�@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     0q@     ȁ@      8@     �K@     @|@     �U@     ��@      m@     @�@     �v@      9@             �R@     �d@      @      @      ^@      @     �z@      E@     pq@      T@      @              H@     �S@      @      @     �P@      @      Z@      ?@     @Z@      G@      @              5@     �A@      @       @      9@      @      H@      4@     �E@      8@       @              @      $@                      @       @      2@      @      &@       @                      1@      9@      @       @      3@      @      >@      0@      @@      6@       @              ;@      F@              @     �D@              L@      &@      O@      6@      �?              "@      4@                      &@              ?@      @      8@      "@      �?              2@      8@              @      >@              9@      @      C@      *@                      :@     @U@      �?       @      K@       @     t@      &@     �e@      A@      �?              �?      ,@      �?              0@       @     �V@      �?      A@      "@                      �?      &@                      "@       @      M@              6@      "@                              @      �?              @              @@      �?      (@                              9@     �Q@               @      C@             �l@      $@     �a@      9@      �?              @       @               @      @             @S@       @      ;@      �?      �?              3@     �O@                     �@@             @c@       @     @\@      8@              &@      i@     Py@      4@      H@     �t@     �S@     P�@     �g@     ��@     �q@      5@      @      K@     �d@       @      ,@     @]@      2@     �u@     �O@     �n@      \@      @      @      0@      ?@      �?              <@      @     �I@      ,@     �E@      <@      @      @      @      *@      �?              8@      �?      4@      *@      .@      5@      @              &@      2@                      @       @      ?@      �?      <@      @              �?      C@     �`@      @      ,@     @V@      .@     �r@     �H@      i@      U@       @              1@     �S@      @      @     �O@      (@     `d@      5@     �`@      K@              �?      5@     �K@      @       @      :@      @     �`@      <@      Q@      >@       @      @     `b@      n@      (@      A@     �j@     �N@     �m@      `@     �q@     �e@      .@       @     �M@      \@      @      3@      S@      3@     �V@     �E@     �[@      N@      &@       @     �@@      O@      @       @      C@      1@      <@      B@      C@     �B@       @              :@      I@      �?      &@      C@       @     �O@      @      R@      7@      @      @      V@      `@       @      .@     `a@      E@     `b@     @U@     �e@      \@      @      @      Q@      Z@      @      ,@     �X@      A@     �P@     �R@     �U@     @S@      @              4@      9@      @      �?      D@       @     @T@      &@      V@     �A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ΕhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��"=M@�	           ��@       	                    �?�����@z           �@                           �?C�=6�@�           8�@                           �?�|��@.           P~@������������������������       ��/�b'@�            �l@������������������������       �,"<�@�             p@                          �<@j8p���@m            @d@������������������������       ��(��A�@f            �b@������������������������       ���^~@             &@
                           @��}��y	@�            �@                          �2@iR/�V	@Z           �@������������������������       ���A�]Q@�            pq@������������������������       ���Iw:�	@�           ��@                          �:@Z��	E	@�            �h@������������������������       �9`�?��@k            �c@������������������������       �`=
6@             D@                          �6@��&��@R           �@                           @4y���@	           �@                           @k�`ۦR@�            �p@������������������������       ���?)DB@�            �i@������������������������       �h޹���@'            �N@                            �?��ò.�@X           ؍@������������������������       �@q30=��?v            �i@������������������������       ��!|h�a@�           h�@                          �>@JF���@I           �@                            @�#پ��@1           `}@������������������������       ���(ڱ@�            �w@������������������������       �HK�8�1@:            �V@                           @Z�	d�@             C@������������������������       ��|�7�S�?             3@������������������������       ��s��Tq@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �q@     ��@      =@     �N@     P|@     �U@     �@     �h@     ��@     Pv@     �A@      8@     @g@      t@      6@      H@     �s@     �Q@     �w@     �c@     Px@     �n@      :@      �?      M@     �S@       @      $@      T@       @     �b@      @@     @c@     �P@      @      �?     �H@      Q@       @      "@     �P@      @     �V@      9@      [@     �K@      @      �?      0@      =@       @      @      ?@      @      H@      0@      H@      :@       @             �@@     �C@              @      B@              E@      "@      N@      =@      @              "@      &@              �?      *@      @      N@      @      G@      &@      �?              "@      &@              �?      &@      @      N@      @      F@      "@                                                       @                      @       @       @      �?      7@      `@      n@      4@      C@     `m@      O@     �l@     �_@     `m@     `f@      3@      0@     �[@     @j@      4@     �B@     �h@      H@     �i@     �Y@     �k@     `c@      .@       @      2@      F@               @      B@             �P@      ;@     �H@      A@              ,@      W@     �d@      4@     �A@     `d@      H@      a@      S@     �e@     @^@      .@      @      2@      ?@              �?      B@      ,@      9@      8@      ,@      8@      @      �?      0@      ;@              �?      <@      ,@      5@      1@      *@      1@      @      @       @      @                       @              @      @      �?      @      �?      �?     �W@     @j@      @      *@     @a@      0@     P�@      D@     p{@      \@      "@             �N@      c@      @      "@     �T@      (@     ��@      &@     0r@      L@      @              :@     �I@      �?              (@       @     �Y@      @      F@      .@      @              ,@     �E@                      (@      @     @U@             �B@      &@                      (@       @      �?                      @      1@      @      @      @      @             �A@     �Y@      @      "@     �Q@      @      {@      @     �n@     �D@      @              @      "@               @      1@      �?     �]@             �F@       @                      >@     @W@      @      @      K@      @     �s@      @     @i@     �@@      @      �?      A@     �L@       @      @     �K@      @      ]@      =@     �b@      L@       @      �?      @@     �K@       @      @      F@      @      ]@      :@     �a@     �F@       @      �?      <@     �I@      �?       @      B@      @     @T@      4@     �]@     �A@       @              @      @      �?       @       @             �A@      @      5@      $@                       @       @                      &@      �?              @       @      &@                               @                       @                      �?      @       @                       @                              @      �?               @       @      "@        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�W�chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@>_�y�`@�	           ��@       	                    �?��E~@�           <�@                            �?^�۔v�@�           ��@                           @Q�3+�l@{            �i@������������������������       ��7Q�p�@?            �Z@������������������������       �L^1�?<            �X@                          �1@r����@(           p|@������������������������       ��(�r71@y            `f@������������������������       ���c	�@�            @q@
                          �1@���m�@�           �@                           �?��ɵ	@�            �v@������������������������       �1f��T @F            �]@������������������������       ��I@�            `n@                           @����2r@           ��@������������������������       �됪�h�@L           �@������������������������       ��ƺnM�@�            s@                           �?��A*�@           �@                          �;@����	@f           0�@                            �?����DJ	@�           ��@������������������������       �*w�d3	@�            �m@������������������������       ��U�/	@/            ~@                           �?��*�@	@�            �n@������������������������       ���,o@9            �W@������������������������       �F�H ��	@c             c@                           @yș�_�@�           А@                           �?_�W@�           �@������������������������       �A�`U?@�            @r@������������������������       ����׳+@�           �@                            �?I���@            �I@������������������������       �7M;ߜ@             @@������������������������       �Ag}����?             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     @r@      �@      >@     �M@      |@     �S@     �@     @k@     ��@     �v@      C@       @     �Y@     �n@      $@      0@      e@      1@     ��@     �V@     �y@     �c@      &@             �@@     @R@              @     �E@      @     r@      .@     �c@     �C@      @              @      >@              �?      $@             �T@       @      N@      (@                      @      3@              �?      "@              5@       @     �C@       @                              &@                      �?             �N@              5@      @                      :@     �E@               @     �@@      @     �i@      *@      X@      ;@      @              @      0@                      3@              V@      @      C@       @       @              5@      ;@               @      ,@      @     �]@      $@      M@      3@      �?       @     �Q@     �e@      $@      *@     @_@      (@     pu@      S@     p@     �]@       @              3@      K@       @      �?      5@      �?      a@      3@     �R@      A@                      .@      .@       @      �?      "@      �?      5@      "@      9@      4@                      @     �C@                      (@             �\@      $@     �H@      ,@               @     �I@     �]@       @      (@      Z@      &@     �i@     �L@     �f@      U@       @       @     �C@     �T@      @      $@     �T@      &@      V@     �I@      Y@      N@       @              (@      B@       @       @      5@             �]@      @     �T@      8@              .@     �g@     �r@      4@     �E@     �q@     �N@     �x@     �_@     �w@     �i@      ;@      ,@     @Y@      d@      ,@      ?@      d@      @@     @Z@     �R@     �`@      _@      0@      @     �Q@     �`@      &@      9@      ^@      5@     @W@     �J@     �[@     �P@      *@              ;@     �C@      @      .@     �E@      @      >@      5@      =@      6@      @      @      F@     @W@       @      $@     @S@      1@     �O@      @@     @T@      F@       @      "@      >@      <@      @      @      D@      &@      (@      5@      9@      M@      @       @      @      (@                      .@      @      @      @      @      @@              �?      7@      0@      @      @      9@      @       @      1@      2@      :@      @      �?      V@     `a@      @      (@      ^@      =@     @r@     �J@     �n@     @T@      &@      �?      S@     @a@       @      (@     @\@      6@     �q@     �E@     @n@     �S@      &@              $@      E@      �?              7@      @     @Y@      "@     �U@      *@              �?     �P@      X@      �?      (@     �V@      0@      g@      A@     `c@     �P@      &@              (@      �?      @              @      @      @      $@       @       @                      @      �?      @                       @      @      "@       @       @                      @                              @      @              �?                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�g�PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@z.���j@�	           ��@       	                   �1@dlF��@e           ��@                          �0@����f�@�           X�@                            @[�!���@~            �g@������������������������       �Q���< @f             c@������������������������       �Ϯ#���@             C@                           @�O��#@           �z@������������������������       �6
���%@�            �r@������������������������       ���H��S@X             `@
                          �4@!Dz
4@�           ��@                           �?��aA��@�           ��@������������������������       �oڌ�r@�            �y@������������������������       ��^ӘD @�           8�@                           @��xK[d@�           ̑@������������������������       �A���&p@�           �@������������������������       �r�kG��@)           `}@                           �?AH�w�/	@?           0�@                          �;@��wg��	@3           `@                           �?�v�B<	@�             l@������������������������       �i~���A
@5            @T@������������������������       ����g��@X            �a@                            @���$ޭ	@�            `q@������������������������       �=�y�@^            �d@������������������������       �i�p�		@H             \@                          @@@-�#[�@            y@                           @D����]@�            0w@������������������������       �� <�!\@�            �p@������������������������       ��g��I@G            @Z@                            �?��~\��@             =@������������������������       �YL��J@             *@������������������������       �Ԉ����?
             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �r@     ��@      C@      L@     �{@     �X@     ؏@     �j@      �@      w@      @@      @     �k@     �|@      8@      F@     t@      L@     ��@     �`@     ؂@      m@      1@      �?      6@      X@      �?      @     �G@       @     q@      5@     �[@      D@                       @     �B@                      5@             �U@      �?      6@      .@                      @      >@                      *@             �S@              1@      $@                      @      @                       @              "@      �?      @      @              �?      ,@     �M@      �?      @      :@       @     @g@      4@     @V@      9@                      @     �F@      �?      �?      *@             @b@      $@      O@      .@              �?      @      ,@              @      *@       @      D@      $@      ;@      $@              @      i@     �v@      7@     �C@      q@      K@     h�@      \@     �~@      h@      1@      @     @W@     �d@      2@      3@     �a@      1@     �v@      O@      o@     @[@      @              @@     �M@              �?      A@      �?     �b@      "@     �Y@      ;@              @     �N@      [@      2@      2@     �Z@      0@     `k@     �J@     @b@     �T@      @       @      [@     @h@      @      4@     �`@     �B@     �o@      I@     `n@     �T@      $@      �?     �S@     �Z@      @      2@     �V@      7@     �[@      F@      `@     �M@      @      �?      =@      V@      �?       @     �E@      ,@     �a@      @     �\@      8@      @      @     �R@     �[@      ,@      (@     @^@      E@     @_@     @T@     �d@      a@      .@      @      I@     @T@      "@       @     �L@     �@@     �E@      M@      L@      V@      ,@              ,@      D@      @      @     �@@      (@      7@      B@      8@      ;@      "@              @      (@       @      @      @      "@      "@      (@       @      &@      @               @      <@      �?              ;@      @      ,@      8@      0@      0@      @      @      B@     �D@      @      @      8@      5@      4@      6@      @@     �N@      @       @      1@      *@      @       @      3@      .@      "@      *@      5@     �G@      @      @      3@      <@       @      @      @      @      &@      "@      &@      ,@      �?              9@      >@      @      @      P@      "@     �T@      7@     @[@      H@      �?              7@      ;@      @      @     �K@      @     @T@      7@      Z@     �E@      �?              3@      .@               @     �D@       @      O@      *@     �R@     �B@      �?              @      (@      @       @      ,@      @      3@      $@      >@      @                       @      @                      "@      @      �?              @      @                      �?      @                       @      @                      �?       @                      �?                              @              �?              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ_��
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �4@,���8@�	           ��@       	                   �1@}B�U�
@�           h�@                           @U$���@�           ��@                           �?f�a��@�            �q@������������������������       ���1���?C            @Z@������������������������       ���kV@k             f@                            �?d�خ���?�            �w@������������������������       ��hΕ=�?�            `k@������������������������       ���o��P�?a            �c@
                           @�RdB@�            �@                           �?UI����@�           ؒ@������������������������       �'���@           @{@������������������������       ��_
��@�           �@������������������������       �;���2�@             2@                           �?�V8�ؖ@           ��@                           �?��#.�	@{            �@                          �<@�_�i"�@�            `q@������������������������       �b�4��@�             m@������������������������       ���S�g@             G@                          �:@TZe
@�           P�@������������������������       �7ɜạ	@<           �@������������������������       ����w�	@�            �m@                          �7@�m7c�E@�           x�@                          �6@N܍�Z�@B           �~@������������������������       �b|��@�            �v@������������������������       ���9S�	@V            �`@                           �?�����q@R           �@������������������������       ��y|!l@�             m@������������������������       ��.續�@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     Ps@     H�@      ;@     �L@     �y@     �T@     T�@     �n@     ��@     pu@      8@       @     �Y@     pp@       @      3@     �d@      1@     @�@     �W@     �w@     �a@      @              ;@     �X@              @      H@       @     �q@      3@     �`@     �C@      �?              1@     �I@              �?     �A@       @     �V@      0@     �G@      6@                      @      &@                      ,@             �I@      �?      8@      �?                      ,@      D@              �?      5@       @     �C@      .@      7@      5@                      $@     �G@              @      *@             �h@      @     �U@      1@      �?              �?      ;@              @      @             �\@      @      I@      *@                      "@      4@                      @             @T@             �B@      @      �?       @     �R@     �d@       @      .@     �]@      .@     �x@      S@      o@     @Y@      @       @     �R@     �d@       @      .@     @]@      ,@     �x@     �R@     �n@     �X@       @       @     �A@     �H@      �?      @     �M@      "@     @X@      J@     �R@     �H@       @              D@     �\@      @       @      M@      @     pr@      6@     @e@      I@                              �?                      �?      �?       @       @      @       @      @      ,@     �i@      t@      3@      C@     �n@     �P@     �v@     �b@     �w@     `i@      1@      *@      `@     �f@      0@      =@      a@     �E@     @[@     @[@     ``@     �\@      *@              C@     �H@      @      @     �B@      �?     �H@      5@     �H@      7@       @             �A@     �G@      @       @      ;@      �?      G@      ,@      E@      *@       @              @       @              @      $@              @      @      @      $@              *@     �V@     �`@      *@      7@     �X@      E@      N@      V@     �T@     �V@      &@      @     �Q@     @Y@      "@      4@     �S@      6@      F@     �J@     �N@     �C@      "@      "@      5@      @@      @      @      5@      4@      0@     �A@      5@      J@       @      �?     �S@     �a@      @      "@     �[@      7@      p@     �D@     �o@     @V@      @              D@      S@       @       @      M@      .@     �a@      &@     �]@      8@      @              6@     �H@       @       @     �H@      *@      [@       @      U@      4@      @              2@      ;@                      "@       @     �A@      @      A@      @              �?      C@      P@      �?      @     �J@       @     @\@      >@     �`@     @P@              �?      1@      7@              @      :@      �?     �I@      "@     @R@      ;@                      5@     �D@      �?      @      ;@      @      O@      5@     �N@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�˺}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�9�^}@�	           ��@       	                    @����p@�           T�@                            @�$�-�@�           P�@                           �?�}d@            {@������������������������       ��6l��@a             c@������������������������       ���6�@�            �q@                           �?���@�            @o@������������������������       �:���\	@{            @i@������������������������       �½ϓl@!             H@
                           @�:o�u@�           X�@                           @�UwV0� @           �y@������������������������       ���͇'@v            �f@������������������������       �g(9�|��?�            �l@                           @���Y�@�            �t@������������������������       ��@y�)� @�            `l@������������������������       ����)n@G            �Z@                          �<@Q�9�jj@!           h�@                          �5@��j=�@]           ֠@                          �4@$я�-@�           ��@������������������������       �Ńe(K@�            0w@������������������������       �3D���@�            �v@                           �?�k֤k@�           0�@������������������������       ���	@�           ��@������������������������       �2#�!�@�           h�@                            �?�А���@�            �t@                           �?�q\I~�@:            @W@������������������������       ��;% ��@             7@������������������������       �,�y���@.            �Q@                          �?@��C@�            �m@������������������������       ��8��@d             e@������������������������       ��8"��@&            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �t@     ��@     �@@      G@     �|@     �W@     ��@     @l@     �@     �v@      =@      @     @V@      g@       @      @     �Z@      8@     0@     �G@     �t@     @^@      @      @      K@      W@      @      @     �U@      2@     �c@      D@     �a@      R@      @      �?     �A@      M@       @      �?      I@      @     �X@      A@     �X@     �E@      @      �?      "@      ?@                      4@      �?      ?@      2@      <@      $@      @              :@      ;@       @      �?      >@      @     �P@      0@     �Q@     �@@      @      @      3@      A@       @      @     �B@      (@      N@      @     �E@      =@              @      1@      <@       @      @     �A@      (@      C@      @     �B@      6@                       @      @                       @              6@      @      @      @                     �A@     @W@      @      �?      4@      @     Pu@      @     �g@     �H@      �?              4@     �N@      @              @      @     �j@       @      T@      3@                      "@      B@                       @      @     @V@       @      <@      $@                      &@      9@      @              @             @_@              J@      "@                      .@      @@              �?      *@             �_@      @     �[@      >@      �?              (@      9@                      @              W@      @      T@      @      �?              @      @              �?      @             �A@      �?      >@      7@              .@     �m@     �w@      9@     �C@     �u@     �Q@     ~@     `f@     p{@     �n@      6@      (@     `i@      u@      8@     �@@     �r@      J@     |@     �b@     �y@     �e@      3@      @      I@     �`@       @      "@     �Y@      1@      f@      A@     �b@      D@      "@      @      9@     @P@      @      @     �J@      @     @Y@      6@      M@      9@      @      �?      9@     @Q@      @      @     �H@      ,@      S@      (@     @W@      .@       @       @      c@     @i@      0@      8@     �h@     �A@      q@     �\@     p@     �`@      $@      @     @R@     �Z@      "@      *@      Y@      :@     @Q@      R@     @U@     @Q@      "@      �?      T@     �W@      @      &@      X@      "@     `i@      E@     �e@      P@      �?      @      B@      F@      �?      @     �J@      2@      @@      ?@      ?@     �Q@      @              @      1@                      0@      *@      @      "@      $@      .@      @              @      @                      @       @                      �?      @                      �?      $@                      "@      &@      @      "@      "@      (@      @      @      @@      ;@      �?      @     �B@      @      :@      6@      5@      L@                      .@      :@      �?      @      6@      @      9@      2@      *@     �D@              @      1@      �?               @      .@      �?      �?      @       @      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJo�ahG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��3�$@�	           ��@       	                    �?�8� �x@l           �@                           �?�=w.T@�           �@                            @�n�&U@�            �s@������������������������       �u3cR�@�            @k@������������������������       �c��b@E            �W@                          �4@�%��c�@           @|@������������������������       �l����@�            v@������������������������       ��o5�Ѕ@9            �X@
                           @��!�N@�           ,�@                            @��Bx�@�           0�@������������������������       �� ��@9           P~@������������������������       ���/� �@Q             `@                           �?�M� �@           (�@������������������������       ��YXFq@           �y@������������������������       ��\$ځ@�            `x@                           @�W�߇@5           �@                           �?����4	@�           X�@                           �?2�X���@�            `q@������������������������       �h��d�@K             _@������������������������       ����Ō�@c            @c@                           �?�!'��	@�            �@������������������������       ��9'�>@�             k@������������������������       ���{�	@z           8�@                           @^��D��@�           X�@                            @���{��@           �{@������������������������       ��Ú��@�            �v@������������������������       ��vW�@1             S@                          �7@�����'@r             f@������������������������       �?��c@"            �G@������������������������       �\��ڹ�@P            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     �@      >@      G@      }@      T@     ��@     �j@     ��@      v@      <@      @     @]@     �r@      &@      5@     �j@      <@     ؆@     @X@     �~@     `c@      *@      @     �O@      \@      "@      @     �\@      0@     `e@      J@      _@     �T@       @              ,@      I@       @             �F@      @      R@      <@     �O@      A@      �?              (@      B@                      9@      �?     �G@      3@     �F@      @@      �?               @      ,@       @              4@      @      9@      "@      2@       @              @     �H@      O@      @      @     @Q@      (@     �X@      8@     �N@     �H@      @      @      A@     �C@      @      @      M@      "@      T@      3@     �E@      G@      @      �?      .@      7@      �?              &@      @      3@      @      2@      @                      K@     @g@       @      .@      Y@      (@     ��@     �F@      w@      R@      @              A@     @W@              @      N@      $@     �i@      =@      a@      C@                      >@     �S@               @      K@      $@     �b@      6@     �Z@      ?@                      @      ,@              @      @             �L@      @      >@      @                      4@     @W@       @      "@      D@       @     v@      0@     �l@      A@      @              @     �H@      �?      "@      8@       @      h@      @     �Z@      2@                      *@      F@      �?              0@              d@      $@     @_@      0@      @      &@     `f@     �n@      3@      9@     @o@      J@     r@     �\@     �t@     �h@      .@      &@     �`@      e@      ,@      3@     �f@     �B@     @]@     �X@     `e@     �a@      .@      �?     �A@     �D@               @     �C@             �F@      2@      N@      A@      @      �?      .@      2@              �?      4@              7@      @      4@      3@                      4@      7@              �?      3@              6@      &@      D@      .@      @      $@     �X@      `@      ,@      1@     �a@     �B@      R@      T@     �[@     @[@      (@              $@      A@      �?      @      B@      @      A@      2@     �B@      ?@      @      $@     @V@     �W@      *@      &@     �Z@      >@      C@      O@     �R@     �S@      "@             �F@     �S@      @      @      Q@      .@     �e@      1@     �c@      L@                      7@     �J@      @      @     �B@      .@     �_@      &@      ^@     �G@                      5@     �I@      @      @      ?@      *@     �V@      $@     @Y@      E@                       @       @               @      @       @     �B@      �?      3@      @                      6@      9@       @              ?@             �F@      @     �B@      "@                      @      1@      �?              @              ,@              @      �?                      3@       @      �?              9@              ?@      @      @@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�xhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @HM��@�	           ��@       	                   �8@ǩ�|��@�           إ@                           @k j���@Y           ��@                           �?.�z�y@b           ��@������������������������       ����Fz�@�            �s@������������������������       �X[5W�#@�           8�@                           �?�ү(@�           ��@������������������������       ���l��� @           �z@������������������������       ��pϕ3@�           ��@
                           @��@�           ��@                           �?Ņ���@�            �w@������������������������       �,����p@C            �Z@������������������������       �r�9��@�             q@                           @�2.T@�            `n@������������������������       ���p�=F@P            @^@������������������������       �*��զ@N            �^@                           @���s�@�           t�@                          �8@�j����@           8�@                          �1@��fS�@r           P�@������������������������       �����M@<            �W@������������������������       ��+��0�@6           �~@                          �<@�����	@�            �k@������������������������       ���g���@W             `@������������������������       ��l^��	@9             W@                           �?��G�c1@�            `s@                          �8@se-�@\            @c@������������������������       ��Asa[@J            �^@������������������������       �%0�a���?             ?@                          �4@�t)�@_            �c@������������������������       �+����?,            �Q@������������������������       �)���H�@3            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     s@     ��@      3@      D@     p}@      S@     |�@     �k@     X�@      u@      :@      *@      k@     �w@      &@      6@     pt@     �K@     8�@     �c@     ��@     �l@      (@      @     `c@     0r@      "@      4@      m@      :@     H�@      Y@     p}@     �a@       @      @      Y@     �^@      @      (@     @a@      .@      i@     @R@      i@      U@       @              F@      <@      �?      �?     �@@       @     @U@      "@     �T@      :@              @      L@     �W@      @      &@     @Z@      *@      ]@      P@     @]@      M@       @             �K@      e@      @       @     �W@      &@      �@      ;@     �p@      L@      @              ,@      M@       @       @      ;@             @l@      @      S@      .@       @             �D@     �[@       @      @      Q@      &@     �q@      4@     `h@     �D@      @      @     �N@      V@       @       @     �W@      =@     �W@      M@     �W@     �V@      @      @     �F@      I@       @             �O@      9@      C@     �D@      E@      P@      @       @      0@      3@                      "@       @      "@      @      4@      6@       @      @      =@      ?@       @              K@      7@      =@     �A@      6@      E@       @              0@      C@               @      ?@      @      L@      1@     �J@      :@                      @      ,@               @      2@      @      ;@      @      <@      2@                      $@      8@                      *@      �?      =@      (@      9@       @              @     @V@     `c@       @      2@      b@      5@      o@     �O@     �n@     �Z@      ,@      @      S@     @`@       @      0@     �]@      4@      `@      N@      b@     @V@      &@             �B@     �X@      @       @     �U@      (@     �Z@      D@     �_@      M@      @              @      .@      �?              @              A@      @      9@      @                     �@@     �T@      @       @     �T@      (@     @R@     �A@     �Y@     �I@      @      @     �C@      @@      �?       @      ?@       @      5@      4@      2@      ?@      @      �?      6@      2@              �?      1@       @      2@      *@      (@      3@      @      @      1@      ,@      �?      @      ,@      @      @      @      @      (@                      *@      9@               @      :@      �?      ^@      @      Y@      1@      @              @      &@              �?      (@      �?      M@              J@      &@      @              @      &@              �?      &@      �?     �D@             �C@      &@      @                                              �?              1@              *@                               @      ,@              �?      ,@              O@      @      H@      @                       @       @                      @              D@              2@                              @      @              �?      &@              6@      @      >@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?45�~�W@�	           ��@       	                     �?ZQ.?7o@
           ̒@                          �6@Ƈh�c�@�            �s@                           �?���S��@�             l@������������������������       �1�-A� @H            �_@������������������������       ��zS_�8@G            �X@                          �8@�����U@>            @W@������������������������       ���>.|@            �D@������������������������       ��GӀ%A@%             J@
                            �?#��Wx�@=           ��@                           @~�|���@�            �u@������������������������       �����])@h            �d@������������������������       �Z66s�&@w            �f@                          �=@��Z��;@^           Ѐ@������������������������       �"˖�|�@P            �@������������������������       �T`:�@             :@                          �1@ U�u�?@�           ,�@                          �0@�����N@�             u@                           @��pS%@?            @W@������������������������       �h荍@%            �M@������������������������       �~��_��?             A@                           @h��M9(@�            `n@������������������������       ����3�@D            �\@������������������������       �����#b�?U             `@                           @Ԫӯ�@�           ��@                            �?(XX_�i@�           0�@������������������������       ���	��S@a           ��@������������������������       ��e�w+T@�            �@                            @g�-Y*	@�            �r@������������������������       �b�?�$�@�             k@������������������������       �����@6            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@      �@      8@     �P@     @|@     �P@     ؏@     �o@     ��@     `x@      =@      �?      X@     �a@              @     @Z@      @     �{@      I@     �o@      Y@       @      �?      .@      A@              �?     �A@      @     �_@      (@     �Q@      3@      �?              "@      ;@              �?      .@              Y@      @     �K@      (@                      �?      @              �?      (@              P@      @      @@      @                       @      5@                      @              B@      �?      7@      @              �?      @      @                      4@      @      ;@      @      .@      @      �?               @      @                      (@              0@       @      @              �?      �?      @      @                       @      @      &@      @      &@      @                     @T@      [@              @     �Q@      @     �s@      C@     �f@     @T@      �?              >@     �G@              �?      9@      @     �\@      0@     �R@      B@                      5@      *@                      (@             �F@      ,@      A@      :@                      "@      A@              �?      *@      @     @Q@       @     �D@      $@                     �I@     �N@              @     �F@             @i@      6@     �Z@     �F@      �?             �G@      N@              �?      D@             �h@      3@     @Z@      D@      �?              @      �?              @      @              @      @       @      @              2@     �i@      w@      8@      N@     �u@      N@      �@     @i@     ��@      r@      ;@      �?      1@     �C@                      6@       @     �`@      1@     �T@      7@                       @      1@                      @             �E@       @      $@      @                       @       @                      @              6@       @       @      @                              "@                       @              5@               @                      �?      "@      6@                      .@       @     �V@      .@      R@      1@              �?      @      "@                      $@       @     �@@      ,@      ;@      (@                       @      *@                      @             �L@      �?     �F@      @              1@     `g@     �t@      8@      N@     Pt@      M@     �{@      g@      |@     �p@      ;@      (@     �b@     �q@      7@      M@     �q@     �H@     �x@     �b@      z@      n@      0@       @     �F@      T@      �?      4@     �O@      0@     �]@     �N@      ]@     �O@      @      $@     �Y@     @i@      6@      C@     �k@     �@@     0q@     �U@     �r@     @f@      $@      @     �C@     �H@      �?       @      E@      "@     �H@     �B@      @@      :@      &@      �?      A@      6@              �?     �@@       @      =@      ?@      9@      8@      "@      @      @      ;@      �?      �?      "@      �?      4@      @      @       @       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@6ը�[@�	           ��@       	                    @�DZ�@n           �@                           �?�����@�           $�@                           �?q���@           `z@������������������������       ���O@(@�            �r@������������������������       �FI�,T�@R            �^@                           �?	�<9�@�           �@������������������������       ��Yxa_�@�            �g@������������������������       �:�+N�@+           @~@
                          �0@͘[�@�           ��@                           @q�u��?L            �^@������������������������       �"�4/���?A            �Z@������������������������       ��������?             0@                           @9�4��}@f           �@������������������������       ��Q!��@�            �l@������������������������       �UL�@�           ��@                           �?�����@K           �@                            �?a�֮�:@�           �@                          �6@��dQ�@�            �h@������������������������       �w�y��� @            �C@������������������������       ��z�i@e             d@                          �?@HNUj@J           ؀@������������������������       �)f4s�@?           H�@������������������������       ���+,��@             2@                           @��] �@�            �@                           �?u��T	@�           ��@������������������������       ���%!�@v             h@������������������������       �l�l�<h	@J           P@                            �?	0��%@�            �r@������������������������       ��r���*@.            @P@������������������������       ����yb@�            @m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     @�@      =@      M@     �{@     �W@     ��@     �i@     ��@     @v@     �A@       @     @\@     `s@      (@      <@      j@      G@     ��@     �T@     `~@     @c@      .@       @     �R@     �d@      "@      5@      c@      @@     �n@      R@     @i@     �Y@      $@      @      =@     �P@      @      @     @P@      2@     @[@      :@      J@     �D@       @      @      9@     �I@       @      @      D@      &@     @R@      2@      A@     �A@       @              @      .@      @      �?      9@      @      B@       @      2@      @              @      G@     @Y@      @      1@      V@      ,@      a@      G@     �b@      O@       @              .@      ?@              �?      .@             �N@      @     �I@      *@              @      ?@     �Q@      @      0@     @R@      ,@     �R@      E@     �X@     �H@       @              C@     �a@      @      @     �K@      ,@     �}@      &@     �q@     �I@      @                      9@                                     �P@              9@      @                              2@                                      P@              8@      �?                              @                                      @              �?      @                      C@     �]@      @      @     �K@      ,@     �y@      &@     0p@     �F@      @              2@      C@                      (@      $@     @T@       @      K@      .@      �?              4@      T@      @      @     �E@      @     pt@      "@     �i@      >@      @      $@     @e@      q@      1@      >@     �m@     �H@     @r@      _@     s@     @i@      4@      @     @S@     @`@      @      $@     @X@      5@     �^@     �@@     �`@      W@      (@              :@      =@       @      �?      :@      @     �F@      "@      A@      .@       @               @       @                      @              4@      �?      @       @                      2@      ;@       @      �?      7@      @      9@       @      ?@      *@       @      @     �I@     @Y@       @      "@     �Q@      1@     �S@      8@     @Y@     @S@      @      �?      F@      Y@       @      "@     @Q@      0@     �S@      8@      Y@     �R@      @      @      @      �?                       @      �?                      �?      @              @     @W@      b@      *@      4@     �a@      <@      e@     �V@     @e@     �[@       @      @      T@      X@      @      3@     �Z@      6@      W@     �R@     �X@     @U@       @      �?      $@      <@      @      @      8@             �C@      (@      C@      =@       @      @     �Q@      Q@      @      *@     �T@      6@     �J@     �O@      N@      L@      @              *@      H@      @      �?      A@      @     @S@      0@      R@      9@                      @      "@      @              @      @      &@       @      1@      "@                      $@     �C@      @      �?      <@      �?     �P@      ,@     �K@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���}hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Y�~�0@�	           ��@       	                    �?P�����@x           �@                            �?����@�           �@                           �?9�xer@�             i@������������������������       �XΚ��@7            @V@������������������������       �"�&g'j@K             \@                          �<@x9q��~@(           �}@������������������������       ���0�@            z@������������������������       �������@#             L@
                          �4@��<u	@�           H�@                           �?+gp��
@|           ��@������������������������       �vFh}l@	           0z@������������������������       �X�k�C7@s            `f@                           @����5�	@R           ��@������������������������       �y���	@�           ��@������������������������       �����@T            �`@                           �?�*)w��@K           X�@                           @i	�� @g           ��@                          �4@z�xy��?�            �w@������������������������       � ��O~�?�            �o@������������������������       �%V�fL�@L            �_@                           �?�� ���@t            �f@������������������������       ��
�O�@H            �^@������������������������       �O8�#k@,             N@                           @��M�@�           ��@                           @�Y�O�@           ȉ@������������������������       �q	IHU�@:           �@������������������������       �Φ5�/~@�            �s@                           @�Vl��@�            �v@������������������������       �
nC�!@�            Pt@������������������������       �5i.��@             D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     �@      :@      M@     �|@     @S@     D�@     �j@     ��@     �u@      <@      5@     �j@      s@      2@     �D@     �s@     �M@     �w@      f@     pw@     �m@      8@      �?     �Q@     �W@      �?       @     �T@      @     �d@      ?@     �b@      P@      @      �?      3@      >@              �?      2@      @     �I@      @     �M@      &@       @      �?      @      &@              �?      "@      @      :@       @      8@      @                      *@      3@                      "@              9@       @     �A@      @       @             �I@     @P@      �?      @      P@             @\@      ;@     @V@     �J@       @             �E@     �M@      �?      @      K@             �Z@      8@     �U@      B@       @               @      @              @      $@              @      @       @      1@              4@      b@      j@      1@     �@@     @m@      K@     �j@      b@     `l@     �e@      4@      @      H@     �R@      @      $@     �X@      @     �]@      G@     �\@      P@      "@      @      E@     �D@      @      @     �R@      @     �S@      @@     �R@     �H@      "@              @     �@@      �?      @      9@       @     �D@      ,@     �C@      .@              0@      X@     �`@      *@      7@     �`@     �G@     �W@     �X@     @\@     �[@      &@       @     �T@     �\@      (@      7@     @^@     �E@     @S@     �P@     @Z@     �X@      "@       @      ,@      4@      �?              ,@      @      1@      @@       @      (@       @             @U@     @n@       @      1@      b@      2@     ��@      C@     Pz@      [@      @              9@     �T@               @      :@      @      r@      "@     �Z@      &@      �?              $@     �J@                      0@      @     �j@       @     @R@      @                      @      =@                      @             �c@             �G@      @                      @      8@                      "@      @     �K@       @      :@      @                      .@      >@               @      $@      @      S@      @     �@@      @      �?              $@      6@               @      @      @      M@      @      0@       @                      @       @                      @              2@      @      1@      @      �?              N@     �c@       @      .@     �]@      &@     `w@      =@     �s@     @X@      @             �E@     @[@       @      @     �Q@      @     `r@      0@     �j@     �O@       @             �@@     �L@       @      �?      I@      @     `d@      *@     @`@     �I@       @              $@      J@              @      5@             ``@      @     @U@      (@                      1@      I@      @      &@      H@      @      T@      *@      Y@      A@      �?              $@     �E@      @      &@     �E@      @     �S@       @     �U@      A@                      @      @                      @               @      @      *@              �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���<@�	           ��@       	                    �?�-�z@e           ��@                          �1@�H��ה@�           ��@                           @p�A���?�            Pq@������������������������       �%�O(<�?�            �l@������������������������       ����DYb@             �G@                           @��s�	@D           �@������������������������       ��3+ň�@�            �s@������������������������       �삾�~
 @            �h@
                           �?����@w           ��@                           �?�I;�@=           @@������������������������       ��>�M�w@p            `e@������������������������       ��&d@�            �t@                           @�>a��s@:           ��@������������������������       ���#�C�@�            Px@������������������������       �z�t[�y@M           �~@                           �?|$y�N�@Z           <�@                          �<@0��6�@1           }@                           �?�Q���@�            pw@������������������������       �R��D��@z            �g@������������������������       ���Т�@{             g@                           �?�1��'@<            �V@������������������������       ������@             E@������������������������       �l</?
�@!             H@                           @�[�n�	@)           ��@                           �?�����	@�           ȉ@������������������������       �>��8�@�            �l@������������������������       ����	@u           ��@                            �?�)�+_o@,           P|@������������������������       �BY�+�@B            �W@������������������������       �N��P_@�            pv@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     ��@      8@     �H@     �@     �U@      �@      j@     P�@     �w@      <@      @     @^@     �r@      @      4@      m@      E@     ��@     �U@     �}@     �c@      "@             �B@     �W@               @     @P@      "@      v@      0@     �d@     �F@      �?              @      ;@              �?      8@              d@       @      I@      @                      @      5@                      .@              b@       @      C@      @                      �?      @              �?      "@              0@              (@       @                      ?@      Q@              �?     �D@      "@     �g@      ,@     �\@     �C@      �?              8@      F@              �?      ?@      "@     �U@      "@     �R@     �@@      �?              @      8@                      $@              Z@      @     �D@      @              @      U@      i@      @      2@     �d@     �@@      w@     �Q@     Ps@     �\@       @      @      K@     @Q@      @       @     @X@      0@     �Q@      D@     �S@      K@      @       @      5@      @@      @      �?      @@      @      6@      3@      0@      0@              @     �@@     �B@              @     @P@      "@      H@      5@      O@      C@      @              >@     �`@       @      $@     �Q@      1@     �r@      ?@     �l@      N@       @              ,@     @R@              @      D@      ,@     �Z@      :@     �T@      <@       @              0@     �M@       @      @      >@      @      h@      @     �b@      @@              "@     `f@     �m@      3@      =@     �q@      F@     @q@     @^@      s@     �k@      3@      �?     �F@      O@      �?      @      N@       @      [@      *@     �Z@     �I@      @      �?     �C@      H@      �?       @     �F@       @      X@      @     �X@      =@       @      �?      <@      <@               @     �A@      �?      :@      @     �F@      1@       @              &@      4@      �?              $@      @     �Q@              K@      (@                      @      ,@              @      .@              (@       @       @      6@      �?              �?       @              @      @               @      @      @      (@                      @      @              �?      (@              @      @      @      $@      �?       @     �`@      f@      2@      7@     �k@      B@      e@      [@     �h@     `e@      0@      @     �W@     �^@      ,@      1@     �a@     �@@      O@     @W@     �Z@     @^@      0@              $@      A@      @      @     �E@      @      :@      9@      ?@      G@       @      @      U@      V@      &@      &@     @X@      >@      B@      Q@     �R@     �R@      ,@      �?      D@     �K@      @      @     �T@      @     �Z@      .@     �V@      I@                      3@      $@                      @      �?      6@      �?      6@      (@              �?      5@     �F@      @      @     �R@       @      U@      ,@     @Q@      C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��m�<@�	           ��@       	                   �<@��+�x�@           �@                            �?ghe@�           L�@                          �8@�tSE@�            �s@������������������������       ��`Z���@�            �p@������������������������       �˗l9�C@            �H@                           �?���@           ��@������������������������       �P^��xw@�            �s@������������������������       ��{>���@T           ��@
                          �?@���3@B             ]@                           @�Z�(��@0            �S@������������������������       ���I�j}@&            @P@������������������������       ��"�v3�?
             *@                          �@@8#�G/@             C@������������������������       �8���N�@	             4@������������������������       ����V��?	             2@                          �4@때m[@�           ��@                            @ƾ�p��@�           ��@                          �1@�IYL�N@            p�@������������������������       � M�Z!$@�            Pq@������������������������       �
$��
_@l           ȁ@                           �?b/���@�            �q@������������������������       �u���k�@j            �c@������������������������       �$1$�K�@N            �_@                          �<@
E�U3	@�           \�@                           @��+��@*           ��@������������������������       ��dꡱ�	@�           `�@������������������������       ���2+�#@7           ~@                          �>@�����(	@�            @m@������������������������       ����="�@R            @a@������������������������       ���ޛ�@A             X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     Ps@     ��@      8@     �J@     �}@     @P@     ��@     `l@     �@     �u@     �A@       @      X@      d@      �?      *@     `a@      @     p{@     �H@     �r@     �S@      @       @     �T@     �b@      �?      @      ]@      @     �z@     �C@     �q@      M@      @       @      .@     �G@                      @@      @      \@      @     �T@      1@                      @     �D@                      :@      �?     �Z@      @      R@      &@               @      "@      @                      @       @      @      �?      &@      @                     �P@     @Y@      �?      @      U@       @     �s@     �A@     �h@     �D@      @             �A@      E@      �?      �?     �I@      �?     @R@      7@     �O@      7@      @              @@     �M@              @     �@@      �?     �n@      (@     �`@      2@                      ,@      (@              @      7@              $@      $@      0@      5@      @              @      &@                      &@              @       @      *@      2@      @              @      @                      "@              @       @      $@      2@      @                      @                       @              @              @                               @      �?              @      (@              @       @      @      @                      @                      @      @              @              @      @                      @      �?               @      "@                       @                              3@     �j@     �w@      7@      D@      u@      N@     ��@     @f@     �@     �p@      <@      @     �O@     �c@       @      "@     @`@      &@     @v@     �N@     �m@     �U@      @             �K@     @]@      @      @     �V@       @     �q@      C@     `f@      N@      @              $@      A@               @      5@             @\@      @     �R@      1@                     �F@     �T@      @       @     @Q@       @     `e@     �@@      Z@     �E@      @      @       @      D@      @      @      D@      @      R@      7@      M@      ;@              @      @      3@      @      @      <@      @      8@      1@      >@      3@                      @      5@                      (@              H@      @      <@       @              ,@     �b@     �k@      .@      ?@      j@     �H@      k@     @]@     �p@     �f@      5@      &@     �]@     �h@      $@      8@     @e@     �D@     �h@     �V@     �m@     �a@      5@      $@     @V@      a@       @      2@     �^@      @@     @R@     �Q@      [@      W@      3@      �?      >@      N@       @      @     �G@      "@     @_@      4@      `@      I@       @      @      ?@      :@      @      @      C@       @      2@      :@      ?@     �D@              @      7@      0@      �?      @      :@      @      @      (@      &@      9@                       @      $@      @              (@      �?      &@      ,@      4@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��9XhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��n�&@�	           ��@       	                    �?BGwV��@�           4�@                          �<@�(-��Y@�           h�@                           �?
Ў�N�@u            �@������������������������       �ˮX���@�            0p@������������������������       �S�aBob@�            t@                          @@@�Ui�E@+            @R@������������������������       �x��a�E@#            �M@������������������������       �M|
:~��?             ,@
                           �? {�@	@�           4�@                           �?�,ޱq�	@�           ��@������������������������       �M̳*�@           �{@������������������������       ��:���	@�           (�@                            �?���Lk@�            �x@������������������������       ��©$�8@M            �`@������������������������       �+���%@�            �p@                           @�rq�@L           ��@                            @f[ sI2@�           L�@                          �4@7��0o�@�           �@������������������������       ���\�� @�           �@������������������������       �����_(@           `z@                          �2@]�)h��?\            �a@������������������������       �x�2 ��?            �F@������������������������       ��1ձ��?=            �W@                           �?��hD�%@Y           ��@                           @+�����@�            �q@������������������������       ��
��@�             k@������������������������       �Xʕ0Z@*            @P@                           @x{���)@�             p@������������������������       ���	�@�             m@������������������������       �+>n�dw@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     ��@      5@     �Q@     �{@     �Q@     (�@      m@     ��@     �u@      7@      .@      m@     pt@      0@     �K@     �t@      K@     `w@     `f@     @w@     �l@      3@             �R@     �T@      @      @     �T@      @      c@     �@@      d@      I@       @              P@     �R@      @      @     �P@      @     `b@      <@     �b@     �A@      �?              ?@      >@      @      @      A@       @     �Q@      3@     �G@      0@      �?             �@@     �F@              �?     �@@       @      S@      "@     �Y@      3@                      $@       @              @      .@              @      @      $@      .@      �?              @      @              @      "@              @      @      $@      .@      �?              @      @                      @              �?                                      .@     �c@     �n@      &@      H@     �n@      I@     �k@     @b@     �j@     �f@      1@      .@      _@      e@      &@      C@     �f@      D@     �a@      ^@      c@     �a@      0@             �@@     �P@       @      5@     @R@      (@     �Q@      E@     @Q@      I@      @      .@     �V@     �Y@      "@      1@     �Z@      <@      R@     �S@     �T@     @W@      *@             �A@     �R@              $@     �P@      $@     �S@      :@      N@     �B@      �?              *@      ;@              @      5@      @     �A@      @      (@      $@      �?              6@      H@              @     �F@      @      F@      4@      H@      ;@                     �Q@     �m@      @      .@     �]@      1@     ��@     �J@     �y@      ]@      @              F@     �b@               @     �R@      "@     (�@      9@     `q@     �Q@      @              E@     �a@               @     @Q@      @     �{@      9@     �l@     �P@       @              1@     @R@               @      7@      @     �s@      0@     @_@      B@                      9@     �P@                      G@      @     �`@      "@     �Z@      ?@       @               @      "@                      @       @     �Q@             �G@      @      �?              �?                                              8@              4@                              �?      "@                      @       @     �G@              ;@      @      �?              :@      V@      @      *@     �F@       @     �a@      <@      a@      G@      �?              *@      J@      @      $@      8@      @     �S@      &@     �P@      3@                      "@      F@      @      @      ,@      �?     �Q@      @      L@       @                      @       @              @      $@      @       @      @      &@      &@                      *@      B@       @      @      5@      @      P@      1@     �Q@      ;@      �?              &@      ?@      �?      @      3@      @      P@      1@     �N@      7@                       @      @      �?               @      �?                      "@      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ-vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�E��o@�	           ��@       	                    @����(@           X�@                          �1@��g@+           d�@                           @��)�@�            `r@������������������������       �Y��d72@�            �k@������������������������       ��j<��@,            @R@                           �?G߲�
�@x           ��@������������������������       ��2���@�            �s@������������������������       �Ő'�O	@�           ��@
                           @6���@�           L�@                           @�?	m @�            0p@������������������������       ��"@I@�            �j@������������������������       ���'�>@             F@                           �?ͻ9,�+@A           ��@������������������������       �ou�)X��?�            Pt@������������������������       ��M��q@o           X�@                           @�P���@~           t�@                           �?����Ԛ	@?           ��@                          �8@sO1��o@�            0p@������������������������       ��7�qd;@5            @V@������������������������       �����
@p            @e@                          �9@4�n{��	@�           x�@������������������������       �� (�+	@�            �r@������������������������       �z�N�\�	@�            0v@                           @4#]�(T@?           X�@                            @]�oL�@�            s@������������������������       ��l��F@�            �o@������������������������       �t���&�?             J@                          �>@�[���@�            @k@������������������������       �Zl``3�@t            �h@������������������������       ����#�@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     0r@     �@     �@@      G@     0{@     @Y@     ��@     �l@     ��@     �v@      B@      (@     `c@     `u@      7@      5@     `l@     �G@     (�@     �Z@     (�@     �i@      ,@      (@     @]@     `f@      *@      (@     @c@      A@     �q@     �W@     @p@     �a@      "@      @      .@     �D@       @              :@       @     �V@      4@     �N@     �@@                      @      <@       @              3@             �R@      *@      J@      :@              @       @      *@                      @       @      1@      @      "@      @              "@     �Y@     @a@      &@      (@      `@      @@     �g@     �R@     �h@      [@      "@             �B@     �B@      �?      �?      ;@      @     �U@      *@     @S@     �@@              "@     @P@     @Y@      $@      &@     @Y@      <@     �Y@     �N@     �^@     �R@      "@              C@     `d@      $@      "@     @R@      *@     �~@      (@     r@     �P@      @              .@     �C@      @              "@      $@     @X@      @     �O@      0@      @               @      =@                      "@       @     �U@      �?     �L@      0@                      @      $@      @                       @      $@      @      @              @              7@      _@      @      "@      P@      @     �x@       @     @l@      I@       @               @      G@               @      *@             �f@      @     �O@      (@      �?              5@     �S@      @      @     �I@      @     �j@      @     `d@      C@      �?       @      a@     �i@      $@      9@      j@      K@      n@     �^@      o@     �c@      6@       @      Y@     �_@      @      3@     �b@      F@     @[@     �Y@     �^@      Z@      4@      �?      =@      ?@      �?      @      D@             �J@      0@      I@      =@      @              @      @      �?      �?      *@             �@@       @      8@      @              �?      7@      9@              @      ;@              4@      ,@      :@      :@      @      @     �Q@      X@      @      ,@     �[@      F@      L@     �U@      R@     �R@      0@             �A@      G@      @      (@      O@      @      :@     �@@      C@      ;@      &@      @      B@      I@      @       @     �H@     �B@      >@      K@      A@      H@      @              B@     �S@      @      @     �L@      $@     ``@      4@     �_@     �J@       @              1@      J@              �?     �B@      @      V@      "@     @S@      3@       @              0@     �I@              �?      >@      �?     @P@      "@      N@      2@       @              �?      �?                      @       @      7@              1@      �?                      3@      :@      @      @      4@      @     �E@      &@      I@      A@                      0@      :@      �?      @      2@      @     �E@      $@      H@      8@                      @               @               @       @              �?       @      $@        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�>�LhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@����m@�	           ��@       	                    �?����@�           �@                           �?���@V           �@                           �?�� �@i             e@������������������������       �h��Ϙ�@.             S@������������������������       ����-i�@;             W@                           �?jZ; e>�?�            �w@������������������������       ����3I(�?�             j@������������������������       �q�~t���?k            `e@
                           @ރu<5@+            �@                          �0@�i�G%@           0{@������������������������       �$G���@             D@������������������������       ����#@�            �x@                           @-�O��@           �z@������������������������       �v�E�9@�            �t@������������������������       �1}��>�@<             X@                           @ OLs@!           ��@                          �<@�` Uf	@�           ��@                          �;@�h�@�(	@           ��@������������������������       �Rf��	@�           h�@������������������������       ����}��@/            @S@                            �?�流�@�            �p@������������������������       ���c���@[            �b@������������������������       ���d���@G            @]@                           @�v�u�@l           ��@                          �=@U����@�           x�@������������������������       ����qE@|           (�@������������������������       �'%��k�@             E@                           @R�\_x�@�            pv@������������������������       �Q�xR��@�            �l@������������������������       �]��}�@K             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     0r@      �@      8@      M@     �}@      T@     P�@     �i@     H�@     `x@     �C@      @     �P@     `f@      @      $@     @`@      ,@     �@      O@     ps@      [@      @              .@     �K@              @      F@       @     `o@      (@     �`@      ;@       @              @      4@              @      7@       @      L@      @     �@@      2@                      @      "@                      (@       @      >@      @      (@      @                      @      &@              @      &@              :@       @      5@      .@                      "@     �A@              �?      5@             `h@      @     �Y@      "@       @              @      6@              �?      ,@             @Z@      @     �K@       @                      @      *@                      @             �V@       @     �G@      @       @      @      J@      _@      @      @     �U@      (@     �p@      I@      f@     @T@      @      @     �A@     �L@      �?      @     �M@      $@     @X@      F@      O@      M@      @              @      .@                      @              $@               @       @              @      >@      E@      �?      @     �J@      $@     �U@      F@      N@      L@      @              1@     �P@      @      @      ;@       @     �d@      @     �\@      7@                      &@      J@       @      @      *@       @     �a@      @     �U@      0@                      @      .@      �?              ,@              9@              <@      @              4@      l@     �v@      4@      H@     �u@     �P@     p~@     �a@      }@     �q@     �@@      1@     �e@     @j@      .@     �D@     �n@     �G@     �g@      ]@     `n@     �g@      ;@      ,@      b@     �e@      .@      >@     �k@      C@     `f@     �T@     �j@     �_@      4@      @     �`@     �d@      .@      =@      j@      A@     �d@      T@     �i@      ]@      4@      @      &@      "@              �?      &@      @      (@       @      "@      &@              @      ?@     �B@              &@      ;@      "@      (@      A@      >@      P@      @              &@      1@              @      $@      @      @      2@      2@     �J@      @      @      4@      4@               @      1@      @      @      0@      (@      &@              @     �H@     `c@      @      @     @Y@      3@     �r@      ;@     �k@     �V@      @      @      8@     �X@       @       @     �Q@      @     @j@      &@     �a@      J@      @      @      4@     �V@       @       @     �J@      @     @j@      $@     �`@     �G@      @              @      @                      1@                      �?       @      @                      9@     �L@      @      @      ?@      (@     �U@      0@     �T@     �C@       @              ,@     �G@      @       @      (@      @     �M@      (@      L@      7@                      &@      $@              @      3@      "@      ;@      @      ;@      0@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��2thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�ѢV�@�	           ��@       	                    �?�LK(��@&           h�@                           �? n�S;�@y           p�@                           �?|��l��@�             o@������������������������       �E�c�4>@5             U@������������������������       ���JT�%@j            �d@                            �?���5�X	@�            Pu@������������������������       �� �sV@=            �W@������������������������       �i �˖	@�            �n@
                          �7@���r�@�           0�@                          �3@��ёMu@	           �@������������������������       �"r��d�@#           `|@������������������������       ���T�M�@�            pw@                           @�Ӻ3@�            �p@������������������������       ��B��C@y            �h@������������������������       �K�ST�@+             R@                            @�sCͩ7@q           ^�@                            �?� �d��@�           ��@                          �5@L>��,I@�           ��@������������������������       ��1�Z�@�           ��@������������������������       �[l�	@V           X�@                          �4@ܠHId@�            �x@������������������������       �qe���@o            �f@������������������������       �z�D@�            �j@                          �:@�=6�)�@�            �@                          �4@N䠱w�@W           ��@������������������������       ��=M~@�            pp@������������������������       ��&Ѷ�@�            �p@                           �?B��W	@D            �\@������������������������       �>��_�@             0@������������������������       ��$��?	@9            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �p@     �@      D@      E@     @@     �R@     ��@      i@     h�@     �w@      >@      @     @W@     �k@      8@      2@      j@     �B@     �}@     @R@     �u@      f@      (@      @     �C@      Z@      1@      @     �U@      7@     �W@      E@     �S@     @V@      "@              3@     �A@      @      �?      G@      @     �I@      .@      F@      9@      @              $@      @                       @              :@       @      :@      @                      "@      <@      @      �?      C@      @      9@      *@      2@      4@      @      @      4@     @Q@      ,@      @      D@      0@     �E@      ;@      A@      P@      @              @      ;@              �?      (@      @      $@      (@      @      ,@       @      @      *@      E@      ,@      @      <@      *@     �@@      .@      ;@      I@      @       @      K@     �]@      @      (@     �^@      ,@     �w@      ?@     �p@      V@      @             �B@     �X@      @      &@     �U@      *@     ps@      5@      h@     �H@       @              3@     �J@      �?       @     �D@              g@      *@     �[@      >@                      2@     �F@      @      "@      G@      *@     �_@       @     �T@      3@       @       @      1@      4@              �?      B@      �?     @Q@      $@     �R@     �C@      �?       @      (@      ,@              �?      4@      �?     �P@      @     �I@      <@                      @      @                      0@              @      @      8@      &@      �?      *@     �e@     �q@      0@      8@     0r@     �B@     ��@     �_@     0@     �i@      2@       @     @Z@     �h@      *@      ,@      h@      :@     �x@     @V@     �w@     �b@      (@      @     �T@     @c@      &@      &@     �`@      3@     0q@      S@     pq@     @_@      &@      �?      :@     @S@      @      @      L@      @     �h@      :@     �e@     �M@      @      @     �L@     @S@      @      @     @S@      0@     �S@      I@     �Z@     �P@       @      �?      6@     �F@       @      @      N@      @     �]@      *@     @X@      9@      �?               @      8@                      *@       @     @T@      @      B@      &@      �?      �?      ,@      5@       @      @     �G@      @      C@      @     �N@      ,@              @      Q@     �U@      @      $@     �X@      &@     �a@      C@     �^@     �K@      @      @     �F@     �Q@      �?      @     �U@      $@     �]@      >@     �\@     �F@      @      @      1@      8@              @      @@      @     �R@      ,@     �Q@      4@       @              <@      G@      �?              K@      @     �F@      0@      F@      9@      �?       @      7@      1@       @      @      (@      �?      5@       @      "@      $@      @              @              �?              @              @                      @               @      4@      1@      �?      @       @      �?      1@       @      "@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�ưԕ3@�	           ��@       	                     @��KC�@�           ��@                          �1@dBQ�@�           �@                           @�r��<�@            �|@������������������������       ��)t���@d            `c@������������������������       ��R<@v @�            0s@                           @��?_t�@�           ȃ@������������������������       �J�d��(@-           P~@������������������������       ���@X            �b@
                           @2�7~�A@�            pv@                           �?����@�            @o@������������������������       �rVG7��@'             P@������������������������       �
/���@u            @g@                           @��e�� @D            @[@������������������������       �����!�?             9@������������������������       �e�� @3             U@                           @�����;@           6�@                          �;@G]�:_	@�           Ȗ@                          �7@{��	@�           �@������������������������       �+����@�           �@������������������������       ��1:�@           |@                          �?@���_	@�             s@������������������������       ���?#Ь@�            �m@������������������������       �p���	@-             Q@                           @/�
bP@m           H�@                           @���R��@�           H�@������������������������       ���V^��@           �z@������������������������       ��\� � @�            �k@                            �?�d��3@�             v@������������������������       �ǃ�A@=            �V@������������������������       ��^���4@�            `p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     �@      8@      N@     p|@     @T@     0�@     @m@     �@     �t@      <@      @     �P@     @h@       @      1@     �a@      ,@     ��@     �R@     @s@     �X@       @              H@     �b@      �?      $@     �W@       @     `z@     �M@     �m@     @P@       @              1@      P@              @     �@@      �?      j@      1@     @W@      7@                      "@      :@                      5@      �?     �G@      &@      =@      &@                       @      C@              @      (@              d@      @      P@      (@                      ?@      U@      �?      @      O@      @     �j@      E@      b@      E@       @              *@     �P@              @     �L@      @      e@      <@     �\@      <@                      2@      1@      �?              @       @      G@      ,@      =@      ,@       @      @      3@      G@      �?      @      G@      @     �[@      0@     �Q@      A@              @      *@      @@      �?      @      C@      @     �O@      .@      D@      @@               @      "@      &@                      *@      �?      &@       @      ,@      �?              �?      @      5@      �?      @      9@      @      J@      *@      :@      ?@                      @      ,@                       @             �G@      �?      ?@       @                       @      @                                      (@              @                              @       @                       @             �A@      �?      :@       @              ,@      m@     �u@      6@     �E@     �s@     �P@     �@     �c@     �~@      m@      :@      *@     �e@      j@      .@     �@@     �j@     �K@      i@     @_@     @m@     �d@      6@      @     �`@     �e@      *@      ;@     `f@      C@      e@      Z@     �h@     �X@      3@      @     @W@     @\@      @      7@      _@      0@     @V@     �G@     �^@      M@      $@             �C@      O@      @      @     �K@      6@     �S@     �L@     �R@     �D@      "@      "@      E@     �@@       @      @      A@      1@     �@@      5@      C@     �P@      @      @      7@      <@       @      @      9@      ,@      <@      0@      >@     �N@       @      @      3@      @              @      "@      @      @      @       @      @      �?      �?      M@     �a@      @      $@     @Y@      (@     �r@      A@     @p@      Q@      @      �?     �A@     @V@               @     �N@      @     �k@      2@     �e@      D@      @      �?      <@      J@              �?     �H@      @     @a@      1@     �Y@      A@      @              @     �B@              �?      (@              U@      �?      R@      @                      7@      K@      @       @      D@      "@     @T@      0@     @U@      <@      �?              @       @      @              @      �?     �A@       @      0@      @                      0@      G@      @       @      A@       @      G@       @     @Q@      6@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���uhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����7@�	           ��@       	                    �?�o#7	@�           \�@                          �<@���jZ(@"           ~@                          �3@q��o_�@�            �z@������������������������       �Z'�/#?@c            �c@������������������������       ����z@�            �p@                          �>@��*�H@#             K@������������������������       �_����@             =@������������������������       �:=I���@             9@
                           �?B�<G�	@�           ؑ@                          �:@���%�y@           �{@������������������������       �'����A@�            �w@������������������������       ����@)            �P@                           @4I�B�-
@�           ؅@������������������������       ��#sW�
@�            �@������������������������       �e�U��@7            �V@                          �4@W])���@�           �@                           �?id�ϱ�@           4�@                           @���ҷ3@           }@������������������������       ��pC�M�?�            @v@������������������������       ��yK�ʽ@F            @[@                           �?©||O�@�           ��@������������������������       ����$G�@�            �v@������������������������       �|��e��@�            �x@                           @���_�@�           ��@                           @?�}�@           p�@������������������������       �QRN���@�            Ps@������������������������       ���l�U@3           �}@                           �?���a�@�            pq@������������������������       ��5.�@R             `@������������������������       �QR��|�@c            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     ؀@      @@     �J@     �|@     �Q@     �@      j@     h�@     �v@      B@      1@     �f@     �l@      6@      A@      n@      F@     �n@      ^@     q@     �g@      :@       @     �M@     @P@      @      @      L@      @     �W@      :@     @[@     �K@      @       @      K@     �M@      @       @      H@      @     @W@      5@     �Y@      B@      @              &@      3@               @      5@      @      C@      $@      D@      *@               @     �E@      D@      @              ;@             �K@      &@      O@      7@      @              @      @               @       @               @      @      @      3@                      @      @                      �?              �?      �?      @      *@                       @                       @      @              �?      @      @      @              .@     @^@     �d@      3@      >@      g@      D@     �b@     �W@     �d@      a@      7@      �?      >@      O@      @      .@     @R@      @     @T@     �A@     �Q@     �M@      @      �?      >@      N@      �?      .@      L@      @     �R@      ;@      O@     �C@      @                       @      @              1@       @      @       @       @      4@              ,@     �V@      Z@      .@      .@      \@     �@@      Q@     �M@     �W@     @S@      1@      $@      V@      V@      .@      .@     �X@      =@      K@     �F@     �V@      P@      (@      @      @      0@                      ,@      @      ,@      ,@      @      *@      @             �]@     @s@      $@      3@     �k@      :@     H�@      V@     ��@     �e@      $@              I@     `c@      @      $@     @U@       @     �@     �B@     s@     @S@      �?              2@      I@               @      9@             �k@      (@     @]@      4@      �?              ,@     �@@                      2@             �f@      @     �W@      (@                      @      1@               @      @              C@      "@      7@       @      �?              @@     @Z@      @       @      N@       @     �q@      9@     �g@     �L@                      2@     �E@       @      @      E@      �?      `@      *@      U@      <@                      ,@      O@      �?       @      2@      �?     �c@      (@      Z@      =@                     @Q@      c@      @      "@      a@      8@     q@     �I@     `m@     �W@      "@              K@     �[@      �?      @     �Y@      .@     �k@      A@     �e@     �L@       @              @@      E@              @      F@      &@     �O@      7@     �L@      @@      �?              6@      Q@      �?      �?      M@      @      d@      &@      ]@      9@      @              .@     �E@      @      @      A@      "@      I@      1@      O@      C@      �?              &@      :@       @      @      2@              9@      @      ;@      &@                      @      1@      @      �?      0@      "@      9@      &@     �A@      ;@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�1�qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�ә��@�	           ��@       	                   �4@?�ۚT�@�           ��@                           @3r��:@*           ��@                           �?�@��@K           8�@������������������������       �Ӷ�s�@t             g@������������������������       ���e�@�            �t@                           �?�.m@�           @�@������������������������       ��Y�6q��?�            Ps@������������������������       �T�(�}#@)           0@
                           �?h���&@�           ��@                           �?G��>�	@p           ��@������������������������       ���b�k�@i            �b@������������������������       �)ZT�)
@           �y@                           �?�>�%Y@$           ��@������������������������       �6����@�             p@������������������������       ��6t �@�           Ѓ@                           @"R��f~@�           ��@                           �?��zՕZ@3           ��@                           �?^�<j?@�            �i@������������������������       �>����* @#             L@������������������������       �����U@`            �b@                          �@@ŋ��^�@�           H�@������������������������       ��Cb�5@�           �@������������������������       �_�z|�X@             (@                          �1@-���ݯ@�            0q@                          �0@����ip�?             F@������������������������       ���'Q"�?	             (@������������������������       ��]籝V�?             @@                          �9@F��o.@�            �l@������������������������       ���l�#@l            �e@������������������������       �}�sP@#            �M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     P�@      6@     �M@     0z@      Q@     x�@      k@     �@     �v@      :@       @     @h@      y@      *@      F@     q@      G@     X�@     �a@     �@     �o@      5@      �?     �M@     �g@      @      "@      V@      @     �~@     �N@     �r@     �\@      @      �?     �@@      R@      @      @      L@      @     @]@      F@     �[@     �Q@      @      �?      "@     �A@               @      6@      @      >@      ;@      @@      6@       @              8@     �B@      @      �?      A@      @     �U@      1@     �S@      H@      �?              :@      ]@      �?      @      @@             �w@      1@     @g@      F@       @               @      ;@                      @             �g@      @     @Q@      "@       @              8@     @V@      �?      @      9@             �g@      *@     @]@     �A@              @     �`@     �j@      "@     �A@      g@      D@     �q@     @T@     �s@     @a@      0@      @      O@     @V@      @      6@     @V@      8@     �Q@     �F@     �S@     �M@      ,@      �?      5@      6@               @      .@             �A@       @      A@      "@      @      @     �D@     �P@      @      4@     �R@      8@     �A@     �B@      F@      I@      &@       @     @R@     �^@      @      *@      X@      0@     �j@      B@     `m@     �S@       @              *@      E@      �?              4@      @     @V@      @      O@      3@               @      N@     @T@       @      *@      S@      $@     @_@      >@     �e@      N@       @       @     �U@     @c@      "@      .@     @b@      6@     0q@     �R@      l@      \@      @       @      S@     �_@      @      *@     �^@      4@     �d@     @Q@      b@     �X@      @      �?      *@     �A@              @      8@      @      I@      $@      E@      4@      @              @      "@                      �?              :@      �?      ,@      �?              �?      "@      :@              @      7@      @      8@      "@      <@      3@      @      @     �O@      W@      @      $@     �X@      ,@      ]@     �M@     �Y@     �S@       @      @      O@      W@      @      $@     @X@      ,@      ]@     �L@     �Y@      S@       @      @      �?               @              �?                       @               @                      $@      ;@       @       @      8@       @     @[@      @      T@      ,@                      @      @                      �?              <@              @                                      �?                                      $@              �?                              @      @                      �?              2@              @                              @      7@       @       @      7@       @     @T@      @     @R@      ,@                      @      5@                      1@       @      N@      @     �L@       @                       @       @       @       @      @              5@       @      0@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �4@�n���0@�	           ��@       	                   �1@��p�5@�           �@                           �?��z=��@�           Ѓ@                           @�����:�?�            �m@������������������������       ��pJ�Y�?z             h@������������������������       ��7Ӥ1� @            �E@                            �?X���@�            �x@������������������������       ��C=�@A             V@������������������������       �ODҁW@�            `s@
                           �?9)�A�3@           �@                          �3@y�h���@�             x@������������������������       ����<x@�            �q@������������������������       ��-�۷�@@             Z@                            �?f8$S@           (�@������������������������       �~>N5�@|            �f@������������������������       �bڳ;�'@�           p�@                           @6�>.j@!           �@                           �?�ʂ+[	@0           ��@                            �?�z���@�            �u@������������������������       ��;��@E            �[@������������������������       ���HC:@�            �m@                           @��� +�	@P           �@������������������������       �	��|	@           �@������������������������       �_φ-y�@J            �_@                           @�+��@�           P�@                          �<@�ePq#;@�           ��@������������������������       �-'��@�           ؄@������������������������       �����S@;            �U@������������������������       ����k�@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �s@     ��@      <@      F@     @|@     @S@     ؏@      i@     ��@     pv@     �B@      @     �Z@     0p@      @      .@     @d@      0@     �@     �R@     y@     `c@      *@       @      =@     @S@      �?      �?      L@      �?      q@      .@      a@      D@      �?              &@      7@                      6@             ``@      �?      E@      @      �?              $@      ,@                      *@             �\@      �?      B@      @                      �?      "@                      "@              1@              @              �?       @      2@      K@      �?      �?      A@      �?     �a@      ,@     �W@     �A@                      @      $@                      @      �?     �F@      @      "@      "@               @      .@      F@      �?      �?      <@             �X@      "@     �U@      :@              @     @S@     �f@      @      ,@     �Z@      .@     w@      N@     �p@     �\@      (@              4@      J@                      >@      �?     �d@      (@     �T@      8@      �?              0@     �C@                      .@      �?      ]@      @      Q@      4@                      @      *@                      .@              H@      @      ,@      @      �?      @     �L@     @`@      @      ,@      S@      ,@     �i@      H@     �f@     �V@      &@              &@      4@                      2@      �?     �M@      7@      >@      *@       @      @      G@     �[@      @      ,@      M@      *@     @b@      9@      c@     �S@      @      *@     �i@     Ps@      5@      =@      r@     �N@     �w@     �_@     �x@     �i@      8@      *@     �b@     �i@      1@      5@     �h@      I@     �c@      [@      i@     `a@      5@      �?     �F@     �G@      @      @     �H@      @     �S@      3@     @R@      8@      �?      �?      $@      4@               @      0@       @      =@      �?      ;@      @                     �A@      ;@      @      �?     �@@       @      I@      2@      G@      5@      �?      (@     �Y@     �c@      *@      2@     �b@      G@     �S@     @V@     �_@     �\@      4@       @     @W@     �_@      &@      2@      `@      B@      Q@     @Q@     �^@     @[@      *@      @      $@      ?@       @              5@      $@      &@      4@      @      @      @              M@      Z@      @       @      W@      &@     @k@      2@     �h@     @P@      @              H@     �Y@       @       @     �U@      "@      k@      1@     �h@     @P@      @             �C@     �V@               @     �P@       @     �h@      0@      g@      J@      @              "@      &@       @              4@      �?      1@      �?      *@      *@                      $@       @       @              @       @       @      �?                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��nw�H@�	           ��@       	                    �?�6����@           $�@                           �?=|(z�$@8           �~@                           �?�ծ��@|             g@������������������������       �!:��	@6            �U@������������������������       �p�J�Y@F            �X@                           �?�X��@�            `s@������������������������       ������@Y             c@������������������������       �����$@c            �c@
                          �=@`[	 ��@�           ؆@                            �?�9�X,@�            �@������������������������       ���fI @x             g@������������������������       ��(��@N           @�@                           @އ��F�@             ;@������������������������       ��	�o�� @             $@������������������������       �)q�"@             1@                           @�c��
@�            �@                          �5@�G<	@�           l�@                          �2@�q�Rg6@�           �@������������������������       ���yoza@�            `s@������������������������       �m#[��`@           �z@                           �?�	%8�	@�           ȉ@������������������������       ���[��7@�             j@������������������������       �9|%V�	@t           @�@                           @�T9�@�           ��@                           �?���V�@�           ��@������������������������       ���N,�@              L@������������������������       ���\,�L@�           ؇@                           �?Ҿ�`�@�             s@������������������������       �PK��@
             3@������������������������       �X����@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     @t@     ��@      =@     �K@     �}@      S@     ��@     @i@     �@     �v@      =@             �T@     �c@      @      ,@     �\@      *@     0{@     �B@      q@      U@      @             �K@      S@      @      $@     �O@      @     �]@      4@     @W@      G@      @              ,@      9@                      7@             �M@      @      E@      *@       @              @      .@                      (@              >@      @      ,@      @                      "@      $@                      &@              =@       @      <@      @       @             �D@     �I@      @      $@      D@      @     �M@      ,@     �I@     �@@      �?              4@      8@      @      "@      6@      @      7@      @      6@      1@                      5@      ;@              �?      2@              B@       @      =@      0@      �?              <@     �T@              @      J@       @     �s@      1@     �f@      C@      @              :@      T@              @     �H@       @     ps@      (@     �f@      ?@      @                      5@              �?      &@      @      T@             �L@      $@                      :@     �M@              @      C@      @     �l@      (@     �^@      5@      @               @       @                      @              @      @      �?      @      �?               @                               @              �?      @                      �?                       @                      �?              @      �?      �?      @              .@      n@     Py@      8@     �D@     pv@     �O@      �@     �d@     x�@     �q@      6@      .@     �d@     �l@      2@      <@     �m@     �K@     �i@     �a@      n@     �i@      3@      @      K@      [@       @      (@     �]@      1@     �`@     �K@     �`@      V@      @      @      >@     �F@      �?      @     �H@       @      Q@      =@      G@     �@@               @      8@     �O@      @      "@     �Q@      .@     @P@      :@     @V@     �K@      @      "@     @\@     �^@      $@      0@     �]@      C@      R@      V@     @Z@     �]@      0@              ,@      7@      �?       @      A@      @      =@      6@      <@      F@       @      "@     �X@     �X@      "@       @      U@      A@     �E@     �P@     @S@     �R@      ,@             �R@     �e@      @      *@     �^@       @     0u@      6@     �q@      S@      @             �F@     �_@      �?      �?     @V@      �?     �q@      1@     �i@      H@      @              @      ,@              �?      @      �?      (@      �?      ,@                              C@      \@      �?             �T@             �p@      0@     �g@      H@      @              =@     �H@      @      (@     �@@      @      L@      @     �T@      <@                      �?      �?                      @      @       @                      @                      <@      H@      @      (@      <@      @      K@      @     �T@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ։�chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�H��c@�	           ��@       	                   �;@
Χ��p	@�           �@                           �?����=�@H           8�@                          �7@8��φ@           �z@������������������������       �,�%Q�@�             t@������������������������       ��q�FB@@             Z@                           @C�>K�	@B            �@������������������������       �	�]ph	@           h�@������������������������       �|!�qL�@�            ps@
                           @ݠ;e
@�            �n@                           �?lD�}{	@u             f@������������������������       ����p>@4             S@������������������������       �u���&�@A            @Y@                          �?@��>��	@,             Q@������������������������       �V����@!            �I@������������������������       ��o���@             1@                          �2@@�Ɲ �@�           �@                           �?ਾ50�@�           Ȇ@                           @l'R$�a�?�            �r@������������������������       ����� @E             [@������������������������       ��]�2��?q             h@                            �?N�S�m@           �z@������������������������       �!�@?            �Z@������������������������       ��̃�n�@�            0t@                          �7@�;��@�           ��@                           @x$��@v           @�@������������������������       ��Og\�@	           Pz@������������������������       �
���.X@m           �@                           @������@n           (�@������������������������       �����@_             a@������������������������       �xr8�?@           �{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     0r@     ��@      >@      H@     �|@      V@     (�@     @k@     ��@     �t@     �E@      3@     `d@     0p@      8@      8@      n@      L@     �h@      b@     �p@     �e@      A@      "@      a@     �k@      1@      ,@      k@      G@      g@     �^@     �m@      _@      <@              C@      S@       @             �L@      @     @U@      8@     �X@      B@      @              8@      H@      �?             �B@      @     �Q@      2@     �U@      @@       @              ,@      <@      �?              4@              .@      @      (@      @      @      "@     �X@      b@      .@      ,@      d@      E@      Y@     �X@     �a@      V@      6@      "@      O@     �Q@      &@      $@     �]@      @@     @R@     �J@      [@     �P@      @             �B@     @R@      @      @     �D@      $@      ;@      G@      @@      6@      .@      $@      :@     �C@      @      $@      8@      $@      ,@      6@      :@     �I@      @       @      7@      B@      @      @      .@      @      $@      (@      1@     �B@      �?       @      @      8@      @      @      @      @      @       @      @      *@              @      2@      (@      @      �?       @      �?      @      $@      &@      8@      �?       @      @      @              @      "@      @      @      $@      "@      ,@      @       @      �?      �?              @       @      @      @      @      "@      &@                       @       @                      �?              �?      @              @      @      �?      `@      u@      @      8@      k@      @@     ��@     @R@     ��@      c@      "@              ;@     @Z@      @      @      C@       @     `t@       @     �e@     �D@      �?              @     �@@                      "@             �d@             �Q@      .@      �?              @      4@                       @             �G@              <@       @                      @      *@                      @             �]@              E@      @      �?              4@      R@      @      @      =@       @      d@       @      Z@      :@                       @      7@              �?       @       @     �J@       @      *@       @                      2@     �H@      @      @      ;@              [@      @     �V@      2@              �?     @Y@     �l@      @      4@     @f@      >@     �{@     @P@     �x@      \@       @              M@     �b@      @       @     �Y@      5@     �s@      <@     �o@     �J@      @              ;@     �P@       @       @     �J@      0@     �X@      5@     �Y@      ;@      @              ?@     �T@      �?      @      I@      @     @k@      @     �b@      :@       @      �?     �E@     �T@              (@     �R@      "@     �^@     �B@     `a@     �M@      �?              (@      4@              @      3@       @      3@      *@      6@      8@              �?      ?@      O@              @      L@      @      Z@      8@     @]@     �A@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ~БBhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �<@ �>?�$@�	           ��@       	                    @�)�2�@�           �@                          �3@��CcN@�           ��@                           @�kgO��@�           ��@������������������������       ��C=�Ew@�           x�@������������������������       ����\a� @             *@                           �?�8��@           ��@������������������������       �Jb�f\	@H           (�@������������������������       �hk"��@�            �s@
                            @Fۼ�@)           8�@                          �4@Q�u�X�@�           �@������������������������       �ݒCk�f@�           H�@������������������������       ��n��8T@�           ��@                          �:@XY����@�             q@������������������������       �Mt��@[@�            0p@������������������������       ���&��?             .@                            �?|��$�	@�            �s@                           @<���8@m             f@                            �?Y����@B            �X@������������������������       �ᡩ��@#             J@������������������������       ��q�w��@            �G@                           �?O@�G@+            @S@������������������������       ��|O4l?@             ,@������������������������       ��NuƄ@#            �O@                           �?�9H,�<
@`            �a@                          �?@�R����@)             O@������������������������       ��'	�F�@             D@������������������������       �_Q!��@             6@                           @YHa4@�	@7            �S@������������������������       �J�`��j@&             K@������������������������       �����@z@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     0r@     ��@      9@      L@     `{@     �R@     ��@     @l@     `�@     Pv@      >@      (@     �p@     �@      2@      E@     �x@     �L@     ��@      g@      �@     Pr@      >@      (@     �g@     Pr@      .@      ?@     Pp@     �A@     Pv@     `b@     �v@     �g@      9@      @     �F@      Z@       @       @     �P@      @      e@     �F@     �b@      P@      @       @     �F@     @Y@       @       @      O@      @      e@     �F@     �b@     �O@       @      �?              @                      @                                      �?      @      "@     �a@     �g@      *@      7@     @h@      <@     �g@     �Y@     �j@     @_@      4@      "@     �[@     �b@      &@      2@     @b@      2@     �_@      S@     �b@      X@      4@              @@     �C@       @      @      H@      $@      O@      :@      P@      =@                     @S@     �k@      @      &@     @a@      6@     ��@     �B@     0{@      Z@      @             �Q@     �h@       @      @     �\@      4@     �@     �A@     0v@     �W@      @             �B@     �X@      �?      @      F@      @     0t@      ,@     �i@     �F@      �?             �@@      Y@      �?      �?     �Q@      0@     �f@      5@     �b@     �H@      @              @      8@      �?      @      7@       @     �]@       @      T@      $@      �?              @      8@      �?              7@       @     @[@       @      T@      $@      �?                                      @                      "@                                      @      :@      <@      @      ,@     �C@      1@      ?@      E@      F@      P@              �?      0@      .@              @      1@      "@      ,@     �@@      :@     �C@                      @      *@              @      "@      @      $@      .@      @      <@                      @      &@               @      @      @       @      @      @       @                       @       @              @       @      @       @       @      @      4@              �?      &@       @                       @      @      @      2@      3@      &@                      @      �?                                      @      @       @                      �?      @      �?                       @      @      �?      .@      1@      &@              @      $@      *@      @       @      6@       @      1@      "@      2@      9@              @       @      @      @      @      $@      @      @              &@      (@                              @      @      �?      @      @      @              @      @              @       @                       @      @                              @      @                       @      @      @      @      (@      @      &@      "@      @      *@                      @      @      @      �?      @      �?      @       @      @      (@                       @      @              @      @      @      @      �?      �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@�U�B1@�	           ��@       	                    @���}2@a           N�@                           �?�3�|�@�           (�@                           �?E2��H@*           `}@������������������������       ��k�x��@�             k@������������������������       ��M{>;@�            �o@                          �3@�]��v@�           А@������������������������       ���/�@           �|@������������������������       �8��0|@�           H�@
                           @�^t��d@�           t�@                           �?�u��r@�           x�@������������������������       �:��&��?�            �t@������������������������       ���0V��@�           8�@                           @����/@           �z@������������������������       ���{���@�            �u@������������������������       �Ԟ�-�@1            �T@                          �;@�p�"g8	@Z           �@                           �?�۾�@>            @                           @v���	@�             p@������������������������       �X �I�@E            @\@������������������������       �P���8	@_             b@                           @!�v,�@�             n@������������������������       �V$[XQl@H            @Z@������������������������       ���P�}b@R            �`@                           @{r��B	@            {@                          �<@��u�m�@�            pr@������������������������       ��mK�'@/            @S@������������������������       ��Vg�t@�            @k@                           �?���Ȣ�@X             a@������������������������       �B��Y|	@5            @T@������������������������       ��x�L��@#             L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �q@     ��@      8@     �K@     �|@      Q@     x�@      l@     0�@     @w@      ;@      "@     �i@     �|@      &@     �B@     �u@     �G@     @�@     �`@     h�@     �l@      $@      "@     �a@     �o@      "@      :@     `n@     �A@     �r@     �W@     �q@     @b@      @              K@      R@       @      @     �K@      @      a@      ,@      Z@      9@                      3@      ?@       @      @      @@      @     �O@      "@     �G@      @                     �A@     �D@                      7@             @R@      @     �L@      3@              "@      V@     �f@      @      5@     �g@      @@     �d@      T@     `f@     @^@      @      @      6@     �P@      @      @     �O@      "@      \@      A@     �T@     �K@      @      @     �P@     �\@      @      0@     @_@      7@      J@      G@     @X@     �P@      @              P@     �i@       @      &@     @Z@      (@     ��@      D@      u@      U@      @              E@     �b@      �?       @      R@      @     �z@      8@     @m@     �I@      �?              "@      I@                      (@      �?     �e@       @     @R@      @                     �@@     �X@      �?       @      N@      @     �o@      6@      d@     �F@      �?              6@      M@      �?      "@     �@@      @      b@      0@      Z@     �@@       @              *@     �H@              @      <@      @     �`@      &@     @T@      1@      �?              "@      "@      �?      @      @              $@      @      7@      0@      �?      $@     @T@     �`@      *@      2@     �\@      5@     �`@     �V@      c@     �a@      1@              A@     @R@      @       @      N@      "@     @S@     �N@     �X@      M@      .@              :@      G@      @      @     �B@      @      5@      F@      =@      ;@      .@              1@      3@              �?      3@              @      0@      6@      $@      @              "@      ;@      @       @      2@      @      1@      <@      @      1@      $@               @      ;@      �?      @      7@      @      L@      1@     @Q@      ?@                      @      .@              �?      (@      @      :@      @      5@      .@                      �?      (@      �?      @      &@              >@      (@      H@      0@              $@     �G@     �N@       @      $@     �K@      (@      M@      >@     �K@      U@       @      @      8@     �G@       @      @     �C@      @      D@      2@     �B@      O@       @      @      @      ,@      @              @       @      0@      @      *@      $@              �?      5@     �@@      @      @      @@      @      8@      .@      8@      J@       @      @      7@      ,@              @      0@      @      2@      (@      2@      6@              @      "@      @              @      "@      @      $@      (@       @      .@                      ,@      "@                      @      �?       @              $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJЬ9=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @Y\�X�H@�	           ��@       	                     @�^���@�           8�@                           �?M0��@u           l�@                           �?����[	@`           ��@������������������������       ��ׇ�}�@�            �s@������������������������       �-�Q�
@�           ��@                           �?&�V��@           �z@������������������������       ���3��@^            `b@������������������������       �i�x�@�            pq@
                           �?��i��@           �@                           �?���]8@�             n@������������������������       ���e���@#             M@������������������������       ���/���@s            �f@                           �?g�+އ	@~           ��@������������������������       ��0����	@/           �}@������������������������       �rGi�3k@O            @]@                           @^�'��@B           ��@                          �4@V#�Y�@�           ܑ@                           �?C߹��-@�           @�@������������������������       �W,�bI'@�            �w@������������������������       �y�5�Z� @�            �r@                           @ �j�[�@<           �|@������������������������       ��UV�S@�            �s@������������������������       � Å� �@e            �b@                           �?��4Qj@U           ��@                           �?w�mE�@z             i@������������������������       �d&��P	@N            �`@������������������������       �,�#&��@,            @Q@                          �6@������@�            �v@������������������������       ���v�@�             k@������������������������       �G A�@X            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Ps@     `�@      @@      O@     �|@      Y@     �@     `h@     8�@     @t@      9@      1@     `k@     �t@      8@      G@     �s@      T@     `w@     @d@     �x@     �j@      5@      @     @`@     �g@      &@     �@@     �h@     �L@     @l@     �X@     �p@     �a@      *@      @     �W@     �`@      &@      :@     �`@     �F@     �`@     �R@      d@      ]@      (@              >@     �G@      �?      @     �G@      @     �P@      "@     �P@     �B@       @      @     @P@     �U@      $@      4@     �U@      E@     @P@     @P@     �W@     �S@      $@             �A@     �L@              @      O@      (@     �W@      9@      [@      9@      �?              (@      (@              �?      *@              I@      @     �H@      @                      7@     �F@              @     �H@      (@      F@      6@     �M@      2@      �?      (@     @V@      b@      *@      *@     �^@      7@     �b@     �O@     @_@      R@       @              3@      D@      �?      @     �@@       @     �P@      1@      E@      .@                      @      (@                      @              4@       @      ,@      �?                      ,@      <@      �?      @      =@       @     �G@      .@      <@      ,@              (@     �Q@      Z@      (@      "@     �V@      5@     @T@      G@     �T@     �L@       @      (@      M@      T@      &@      "@     �T@      2@     �H@      A@     �Q@      F@       @              (@      8@      �?               @      @      @@      (@      (@      *@              �?     �V@     �k@       @      0@     �a@      4@     X�@     �@@     �y@     �[@      @      �?     �N@     �c@      @       @      S@      ,@     `}@      1@     0q@     @P@      @              ;@     �V@      �?      �?      9@      @      t@      $@     �d@      B@                      2@      C@              �?      3@             `g@       @      U@      :@                      "@      J@      �?              @      @     �`@       @     @T@      $@              �?      A@     �P@       @      �?     �I@      "@     �b@      @     �[@      =@      @      �?      $@     �G@              �?      =@      @     �\@      @     �T@      2@                      8@      3@       @              6@       @      B@      @      ;@      &@      @              =@     @P@      @      ,@     @P@      @     �f@      0@     @a@      G@      �?              @      ?@       @      �?      "@             �V@      @     �F@      .@                      @      5@              �?       @              O@      �?      <@       @                              $@       @              �?              =@      @      1@      @                      :@      A@      @      *@      L@      @     �V@      (@     @W@      ?@      �?              $@      4@       @      @      5@      �?     @Q@       @      Q@      1@      �?              0@      ,@      �?       @     �A@      @      5@      $@      9@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJbhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�s�01@�	           ��@       	                    �?Ͱ�^��@_           Ҡ@                          �:@��u�	@�           ��@                           �?FO�)�@3           ؓ@������������������������       �X���7@�            �x@������������������������       ����:	@4           h�@                            @7�%�%
@�            Ps@������������������������       �G$�3��@t            �f@������������������������       ��İJ�
@L             `@
                          �=@A�K��@l           ��@                            �?i�L���@Y           ��@������������������������       �7<gU�@�            �s@������������������������       �@���"�@�            �l@                           �?���r�@             ?@������������������������       �[�����?             ,@������������������������       �	�O�@             1@                            �?W��[@P           ��@                          �7@m¡�@R           P�@                           @�1�?�@�           �@������������������������       ��"Kd�@P           ��@������������������������       ��C넹�@�            �i@                          �:@��N�!{@z             i@������������������������       ���y��@<            �X@������������������������       �gz��>/@>            �Y@                           �?�h�ݶ�@�           ��@                            @�c#B @�            pr@������������������������       ���Qۧ� @u            �f@������������������������       �}Fe|t��?B            �\@                           @�G��	p@G           x�@������������������������       ��iRjh�@�            �o@������������������������       �`�h�/�@�            0q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     `r@     �@      9@      F@     p|@     �S@     �@     �l@     Ȉ@     pt@     �B@      4@     �j@     �t@      0@      <@     �s@      L@     w@     �g@      w@     �j@      ?@      4@      e@     `n@      .@      7@     �m@      G@     @m@      a@     @p@      e@      :@       @      a@     `i@      "@      1@     �h@     �A@     �i@     �X@      l@     �\@      5@             �B@     �P@      �?      @     �G@       @     �T@      4@     �X@      @@      @       @      Y@      a@       @      ,@     �b@     �@@      _@     �S@     �_@     �T@      2@      (@      ?@      D@      @      @     �E@      &@      ;@     �C@     �A@      K@      @      @      ,@      5@      �?              ;@      @      5@      2@      9@      C@      @      @      1@      3@      @      @      0@      @      @      5@      $@      0@       @             �F@      W@      �?      @      S@      $@     �`@     �I@      [@      G@      @              E@     �U@      �?      @     �R@      @     @`@     �E@     �Z@      G@      @              =@     �L@      �?      @     �B@      @     @Q@      7@     �Q@      ,@      @              *@      =@                      C@      �?     �N@      4@     �A@      @@                      @      @              �?      �?      @      @       @       @               @                       @              �?                      �?       @                       @              @      @                      �?      @      @               @                      �?     @T@     �n@      "@      0@     �a@      7@     ��@     �D@     �z@     @\@      @             �B@      a@      @       @     �O@      ,@     Pt@      9@     �o@     �Q@                      9@      [@      @      @      G@      &@     `r@      $@     �f@     �I@                      0@     �S@      �?              6@      @     �l@       @      a@     �A@                      "@      >@      @      @      8@      @     @P@       @     �F@      0@                      (@      =@              @      1@      @      ?@      .@     �Q@      4@                      @      @              @      ,@      @      2@      $@     �@@      "@                       @      8@                      @              *@      @      C@      &@              �?      F@     �Z@      @       @     @S@      "@      u@      0@     �e@      E@      @              *@      @@                      .@      �?     �d@      "@      K@      @      �?              @      8@                      @      �?      X@      "@      @@      @      �?              @       @                      "@              Q@              6@       @              �?      ?@     �R@      @       @      O@       @     �e@      @     �]@      B@      @      �?      @      A@              �?      C@      @     @U@      @     @P@      $@      @              :@     �D@      @      @      8@      @     �U@       @     �J@      :@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�w�ahG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?u
RD@�	           ��@       	                    @>��ύ,	@�           ��@                          �1@��229�@�           ��@                           @2�~3��@e            `c@������������������������       ��΀8�6@:            �U@������������������������       �H�Cq�@+            @Q@                           �?x�м;	@B           D�@������������������������       �x��6]@&           `}@������������������������       �ę���	@           ؉@
                           @"���@T             b@                          �7@gFF�@B            @]@������������������������       ��*�M�@*            �R@������������������������       ��ue)�@             E@                           �?�uׅ�d@             <@������������������������       �V@���@             *@������������������������       � �ܤ�@
             .@                           �?�[�ګ@�           �@                          �4@\&�A@�           ��@                           @�T6����?           P}@������������������������       �m��>�@;             Y@������������������������       �xEp���?�            w@                            @:S�J��@�            t@������������������������       ���[�(�@�            `o@������������������������       ����̳��?(            �Q@                           �?Έ2�H�@�           ؗ@                           @;���}@>             Z@������������������������       �)��갦@0            @S@������������������������       �0/�jsx @             ;@                           �?|B	Ӻ@�           8�@������������������������       ���tM64@�           ��@������������������������       �8�a�"@�           ȇ@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@      r@     Ѐ@      <@      M@     �{@     @Q@     ��@     �h@     ؊@     �v@     �B@      ,@     �d@      n@      2@     �A@     @m@     �B@     @l@     �`@     �p@      h@      @@       @     @c@     �j@      2@     �@@     �j@      A@      k@     �Z@     pp@     �d@      :@      �?      @      =@               @      =@              B@      @      A@      1@                      @      0@                      2@              7@      @      0@      @              �?              *@               @      &@              *@              2@      &@              @     �b@     @g@      2@      ?@     �f@      A@     �f@      Z@     �l@     �b@      :@       @      C@      U@      �?       @      N@      @     �X@      <@      V@     �J@      @      @      \@     �Y@      1@      7@     �^@      =@     @T@      S@     �a@      X@      6@      @      &@      :@               @      6@      @      $@      9@       @      :@      @       @       @      :@               @      2@      @       @      4@      @      7@      �?              @      5@               @      0@       @      @      @       @      0@               @       @      @                       @      �?       @      0@      @      @      �?      @      @                              @               @      @       @      @      @       @                                      �?                      @              @      @       @      @                              @               @      �?       @               @             �^@     �r@      $@      7@     `j@      @@     ��@     �P@     `�@     �e@      @              <@      V@              @     �I@      @     pw@       @      i@      <@      �?              0@      G@              @      7@             `n@      @      ^@      *@      �?              @      $@                      $@              @@              B@      @                      "@      B@              @      *@             `j@      @      U@       @      �?              (@      E@                      <@      @     �`@      @      T@      .@                      &@      D@                      5@      @     @X@       @      N@      *@                      �?       @                      @             �A@      @      4@       @                     �W@      j@      $@      3@      d@      9@     �y@     �M@     @x@     @b@      @              "@      ,@              @      0@      @      $@      $@      ;@      &@                       @      ,@              @      @      @      $@      @      3@      @                      �?                              "@                      @       @      @                     �U@     `h@      $@      0@      b@      5@     y@     �H@     �v@     �`@      @             �B@      X@      @      (@     �T@      @      d@      8@     �d@      Q@      @             �H@     �X@      @      @     �N@      ,@      n@      9@     `h@     �P@      �?�t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJaz�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?~�|r@�	           ��@       	                   �4@N�=`Pp	@            `�@                            �?THjK�F@v           ��@                           �?+�*$o@b            �b@������������������������       ���:?V@!            �H@������������������������       ��9�h@A            �X@                           @�䂨Q�@           �{@������������������������       �1�p���@�            `u@������������������������       ���Xu	@=             Z@
                           �?mU�o��	@�           �@                           �?'�R�b�@�            �q@������������������������       ��r��v�@F            �[@������������������������       �(�
�ƭ@m            �e@                           �?nDj]�
@�           H�@������������������������       �X�B紪	@�            @p@������������������������       � �;ҽ
@7           P~@                           @���@�           �@                            @��Q��@o           �@                            �?������@           �x@������������������������       ���1�@k             d@������������������������       �6�^�#@�            �m@                          �6@w��%C�@h            �e@������������������������       ��"9V�t@<             Z@������������������������       �<O�g@,            �Q@                           @m�8w^H@S           К@                          �2@Mrg�3@�            �@������������������������       ��T?Ǽ @           z@������������������������       �t��(@�           8�@                            @ivSg��@W           `�@������������������������       ��D+_�@           �z@������������������������       ������@P            ``@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �s@     ��@     �A@     �G@     P|@     �U@     p�@      l@     @�@     `w@      <@      7@     `e@     �m@      6@     �@@     �n@     �I@     `l@      a@     `o@     `i@      8@      $@      I@     �T@      @      @     �S@       @     �^@      F@     @[@     �Q@       @              "@      7@                      2@      �?      E@      *@      8@      *@      @              �?      $@                      @              2@      @      (@       @                       @      *@                      .@      �?      8@      $@      (@      &@      @      $@     �D@      N@      @      @     �N@      @      T@      ?@     @U@     �L@      @      @      @@     �A@      @      @      I@      @     @R@      .@     @R@      F@              @      "@      9@      �?      �?      &@      @      @      0@      (@      *@      @      *@     @^@     `c@      .@      =@     �d@     �E@     @Z@     @W@     �a@     �`@      0@      �?      ?@     �E@      �?      $@      G@      �?     �B@      *@      O@     �B@      @      �?      ,@      *@                      5@              :@       @      5@      &@      �?              1@      >@      �?      $@      9@      �?      &@      &@     �D@      :@       @      (@     �V@      \@      ,@      3@     �]@      E@      Q@      T@      T@      X@      *@      @     �A@      F@      @      @      D@      ,@      .@      >@      2@     �E@      @      "@     �K@      Q@      @      *@     �S@      <@     �J@      I@      O@     �J@       @      �?     `b@      s@      *@      ,@      j@     �A@     X�@     �U@     h�@     `e@      @              F@      W@       @      @     @P@      $@     @a@     �F@     �^@     �G@       @              C@     �O@              @      L@       @     @U@      <@     @W@      5@       @              @     �@@              �?      2@       @     �C@      &@     �@@      .@       @              @@      >@              @      C@      @      G@      1@      N@      @                      @      =@       @      �?      "@       @     �J@      1@      >@      :@                      �?      *@       @      �?      @       @     �B@      &@      8@      $@                      @      0@                      @              0@      @      @      0@              �?     �Y@     �j@      &@      "@      b@      9@     �@      E@      y@      _@       @      �?      Q@     �a@       @       @     �W@      0@     �}@      .@     `p@     �S@       @              .@      L@      �?              .@      �?     `j@      @     �T@      =@              �?     �J@      U@      �?       @      T@      .@     �p@      "@     `f@     �H@       @             �A@      R@      "@      @     �H@      "@     @d@      ;@     �a@      G@                      @@     �O@       @      @      C@       @      [@      9@     �Z@      @@                      @      "@      �?       @      &@      �?      K@       @      A@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ ��
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@'R�;�;@�	           ��@       	                    @���t�@�           ��@                          �1@|LE�&�@1           �~@                           @�Ȱ�[@�            q@������������������������       �h�g�@Q            �`@������������������������       ���@Z            �a@                           �?��e�@�            @k@������������������������       �I�"m�@3            �U@������������������������       �J�e���@S            ``@
                            �?c�|.U� @a           ��@                           @@�}Pf� @�            �t@������������������������       �	Pc�3��?�            `o@������������������������       �q	Ҋ�b@4            �S@                            @g@q] @�            @n@������������������������       �ߤ��l@[            �b@������������������������       �h۪���?9             W@                           �?b�x �@           D�@                          �:@�fu��p	@-           |�@                           �?p��W'Y	@i           @�@������������������������       �A�,@ o@�            �w@������������������������       ��n��	@�           ��@                           @H��X�@�            ps@������������������������       ��<���@�            �p@������������������������       ��d��5�@            �D@                           �?�~^=��@�           �@                           @3{�Cl�@*           �|@������������������������       ��Zx%k�@            �g@������������������������       �"�Ej�` @�            �p@                           @	�&��@�           �@������������������������       � ����~@�            �q@������������������������       ��89�@�           �@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     s@     ��@      3@     �F@     0}@     @U@     ,�@     �l@     `�@     Py@      ?@       @      D@     �\@               @     �[@       @     0{@      I@      l@     �Q@      @       @      :@      J@              �?     @T@       @     �a@     �E@     @Y@      C@      @              .@      ;@              �?     �@@             �W@      :@      M@      2@                      @      @                      (@             �F@      3@      ?@      (@                      "@      4@              �?      5@              I@      @      ;@      @               @      &@      9@                      H@       @      G@      1@     �E@      4@      @       @      @      @                      :@              8@      @      ,@      @       @              @      2@                      6@       @      6@      *@      =@      0@       @              ,@     �O@              @      =@             `r@      @      _@      @@       @              @     �A@              @      .@             @e@       @     @Q@      :@                      @      ;@                      @             @b@       @     �H@      0@                               @              @      $@              8@              4@      $@                       @      <@                      ,@              _@      @     �K@      @       @              @      5@                      @              S@      @      =@      @       @              @      @                      @              H@              :@      �?              ,@     �p@     �y@      3@     �B@     Pv@     �T@     ��@     `f@     X�@     �t@      9@      ,@     �e@     `f@      *@      6@     �g@      M@     `c@     �^@     �e@      h@      3@      @     @_@     �b@      $@      4@      b@     �C@      `@     �W@     �b@     �]@      1@              >@     �O@      �?      "@      M@      @     @Q@      9@     �Q@     �E@      �?      @     �W@     �U@      "@      &@     �U@     �@@     �M@     �Q@     @S@      S@      0@       @     �H@      >@      @       @     �F@      3@      ;@      <@      8@     �R@       @       @     �G@      :@      @       @     �D@      1@      9@      0@      8@     �P@              @       @      @                      @       @       @      (@              @       @             �V@     @m@      @      .@      e@      9@     �{@      L@     �u@     �a@      @              1@     �S@               @      >@      @     �e@      $@      _@      .@      �?              .@     �A@                      2@      @     �I@      @     �J@      @      �?               @     �E@               @      (@      �?     @^@      @     �Q@      "@                     �R@     �c@      @      *@     @a@      2@     q@      G@     `l@     �_@      @              1@      J@              @     �F@      @     �D@      9@     �J@      A@      �?             �L@      Z@      @      @     @W@      (@      m@      5@     �e@     @W@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�y�Ӱ[@�	           ��@       	                   �:@� �E	@�           |�@                           �?�bh@�@4           ��@                           �?��&/��@E           P�@������������������������       �ڎ%a#a@c            �c@������������������������       ���I��@�            �v@                           @ڣ�U��	@�           �@������������������������       ������!	@w           ��@������������������������       �����	@x            `h@
                           @Qhݫ�@�            @s@                           �?�ϭ+@�            @q@������������������������       �u��u@>            �V@������������������������       �;��ǋU@v            @g@                          �<@1�0�@             @@������������������������       �|R��>�?             0@������������������������       �|R��>@
             0@                            �?�]jOZM@�           ԡ@                           �?㕐�_@[           h�@                          �8@�Z� *@s            `e@������������������������       ��6�*��?f             b@������������������������       �Vh�^�@             ;@                           @�v��@�             v@������������������������       ��t^=�0@�             u@������������������������       �����@	             0@                          �8@ĿԾ�P@j           t�@                           @)*���@�           ��@������������������������       ������@�            �t@������������������������       ����)ծ@�           Đ@                            �?�2�N��@�            �u@������������������������       ���<B�?@I             ^@������������������������       ��P�
@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     ��@      <@      N@     �}@     �V@     `�@     `k@     ��@      v@      @@      *@     `d@     �k@      2@     �@@      q@     �J@      n@     �_@     �p@     �h@      7@       @     @a@     @g@      ,@      ;@     @j@      @@     @l@     �Y@      m@     �_@      5@              B@     �T@      �?      "@      T@      @     @^@      ?@      [@     �E@      @               @      9@                      1@              H@      @     �F@      "@                      <@      M@      �?      "@     �O@      @     @R@      :@     �O@      A@      @       @     �Y@     �Y@      *@      2@     @`@      :@     @Z@     �Q@     @_@     �T@      1@      @     �S@     @Q@      "@      $@     �Z@      7@     �T@      E@     �X@     �R@      @      �?      8@      A@      @       @      7@      @      7@      =@      :@      "@      &@      @      9@      A@      @      @      O@      5@      .@      9@      B@     @R@       @      @      8@      ?@      @      @     �L@      2@      *@      *@      A@     �Q@       @       @      @      @       @              9@      �?      @       @      2@      8@      �?      �?      1@      ;@       @      @      @@      1@      "@      &@      0@     �G@      �?       @      �?      @                      @      @       @      (@       @       @                                                      @               @       @      �?       @               @      �?      @                       @      @              @      �?                      �?     `a@     �s@      $@      ;@     �i@     �B@     ؇@      W@     ��@     `c@      "@              :@     �R@      @      @     �D@      @     @i@      :@     @X@     �C@      @               @      1@      @      �?      @      @      V@             �B@      (@      @               @      1@      @      �?      @      �?     �S@              @@      @                                                               @      "@              @       @      @              8@     �L@       @      @      B@      @     �\@      :@      N@      ;@                      6@      K@               @      B@      @     @\@      7@      N@      8@                       @      @       @       @                      �?      @              @              �?     @\@      n@      @      6@     �d@      >@     ��@     �P@     {@      ]@      @      �?      R@     �j@      @      (@     �\@      :@     �~@     �E@     v@      R@      @              5@     �O@              @     �C@      @      V@      ;@     @P@      3@              �?     �I@     �b@      @      @     �R@      5@      y@      0@      r@     �J@      @             �D@      :@              $@      I@      @     @R@      7@      T@      F@                      5@      *@              @      ,@      �?      (@      $@      <@      0@                      4@      *@              @      B@      @     �N@      *@      J@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJʪhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?UnG��f@�	           ��@       	                    �?Z��w@/           H�@                          �;@Z��+S?@G            �@                           �?�����@            p|@������������������������       �$:9�@�             i@������������������������       �������@�            �o@                           �?\��@'            �L@������������������������       ��&��b@             9@������������������������       ��4u��@             @@
                          �=@)d�@s@�           ��@                          �8@����@�           ��@������������������������       ��ϣ�q @�           ��@������������������������       �������@A            @Z@                          �?@���G��@             4@������������������������       ���T�_ @             $@������������������������       ��	�o�� @             $@                            �?���vc@�           n�@                           @���5a@�           @�@                           �?��'�X;	@!           �|@������������������������       �xl�3@M             _@������������������������       ���'Գ	@�            �t@                           @^�[;�@�            �o@������������������������       �|�ehA�@x            @e@������������������������       �<fw�@3             U@                          �5@�CjZ�D@�           ��@                          �1@��%�k�@�           ��@������������������������       �1��j@�            �l@������������������������       �V�>ӝ@�           x�@                           @�ٹX�	@;           Ћ@������������������������       ��ls4Z}	@]           �@������������������������       �Pّ�@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `s@     `�@     �D@      H@     �{@     �S@     h�@     �i@     p�@     0v@      D@      �?     �W@      h@      @      (@      W@      $@     P~@     �G@     �p@     @V@      @      �?      N@     @W@      �?      $@      O@      @     �Z@      @@     �V@      H@       @              L@     �T@      �?      @     �K@       @      Z@      =@      U@     �@@       @              5@      @@      �?      @      <@       @      J@      3@      <@      (@                     �A@     �I@                      ;@              J@      $@      L@      5@       @      �?      @      $@              @      @      @      @      @      @      .@              �?              @              @      @      @              �?      @      @                      @      @              �?      @              @       @       @      "@                      A@      Y@       @       @      >@      @     �w@      .@     @f@     �D@      �?              A@      Y@       @       @      <@      @     Pw@       @      f@      C@                     �@@      S@       @       @      7@       @     @u@      @     �b@      =@                      �?      8@                      @      @     �@@       @      <@      "@                                                       @              @      @       @      @      �?                                                              @      @      �?      �?      �?                                               @              �?      @      �?       @              1@      k@     �x@      C@      B@     �u@     @Q@     @�@     �c@     �@     �p@     �B@             @Q@     �Y@      @      &@     �V@      0@     �b@      O@     @]@     �R@      1@              I@     @Q@      @      "@      R@      .@      N@      J@      N@     �I@      1@              @      0@              @      8@       @      8@      *@      7@      *@      �?             �F@     �J@      @      @      H@      *@      B@     �C@     �B@      C@      0@              3@     �@@       @       @      3@      �?      V@      $@     �L@      7@                      &@      8@       @              *@             @Q@      @     �C@       @                       @      "@               @      @      �?      3@      @      2@      .@              1@     `b@     Pr@     �@@      9@      p@     �J@     @w@     @X@     �x@      h@      4@      @      K@     �e@      2@      .@      \@      3@     �o@     �D@     `m@     �S@       @       @      ,@      B@       @              ,@             @U@      @      M@      ,@              @      D@     @a@      0@      .@     �X@      3@      e@      B@      f@     @P@       @      (@     @W@     �]@      .@      $@     @b@      A@     �]@      L@      d@     @\@      (@      "@     �R@     �S@      "@      @     @W@      =@      D@     �G@     @S@     �Q@      @      @      3@     �D@      @      @     �J@      @     �S@      "@      U@      E@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�#3&hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�ny,7@�	           ��@       	                    �?]+��E�@|           8�@                           �?�4��$@�           ��@                           @�SCz@�            0v@������������������������       ���Q*@v            �g@������������������������       �û�s��?m            �d@                            �?�XcX� @�            �r@������������������������       ���d��?6            �W@������������������������       ����h:@�             j@
                           @X�{`Fb@�           ��@                           �?a���@r           �@������������������������       �*o����@�            �x@������������������������       ���<�7@u            @g@                           @�[�9��@h           ؁@������������������������       �wf�	�@�            �o@������������������������       ��QK�)N@�            �s@                           �?>�߈a�@/           v�@                          �:@S�P��	@~           ��@                           �?���@�           �@������������������������       �`�H5�@x            �g@������������������������       �$`��Q.	@1           0~@                           @�U�/�	@�            �u@������������������������       ��G��	@�            �m@������������������������       �Ym��"@=            �Z@                           @��OL�@�           ��@                           @+��
H@�           `�@������������������������       ����5R@            �{@������������������������       ���V&Og@y           Ȃ@                           !@���@            �C@������������������������       ��� ��@             3@������������������������       ��4F@             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     ��@      =@      N@      |@      U@     \�@      j@     �@     w@      :@      @     �R@     �j@      @      5@     @g@      2@     ��@     �T@     �x@      `@      @              8@      N@              @     �G@             �t@      *@     �a@      ?@      �?              "@     �A@              @      ;@              f@      $@      R@      3@                      @      7@              @      4@             �Q@       @      D@      0@                       @      (@               @      @             �Z@       @      @@      @                      .@      9@              �?      4@             @c@      @     �Q@      (@      �?              @      (@                                      L@              2@      @                      (@      *@              �?      4@             �X@      @     �J@      @      �?      @     �I@     `c@      @      ,@     `a@      2@     �t@     @Q@      p@     @X@      @      @      B@     @V@      @      $@      W@      .@     �W@     @P@     �X@      N@      @      @     �@@      G@      �?       @     @S@      *@      J@      D@     �P@      F@      @              @     �E@      @       @      .@       @     �E@      9@      @@      0@                      .@     �P@      �?      @     �G@      @     �m@      @     �c@     �B@                      @      D@                      3@      @      V@      @      T@      .@                      (@      :@      �?      @      <@             �b@             �S@      6@              .@     `j@     �s@      6@     �C@     �p@     �P@     x@     �_@     0y@      n@      3@      ,@     �`@     �d@      *@      9@     �a@     �B@     �[@     �S@     @a@     �b@      .@      @     @Y@     �\@      @      *@     �Y@      2@      V@     �E@     �Y@     �Q@      &@              A@      >@       @      @      7@             �D@      @      E@      $@              @     �P@     @U@      @      $@      T@      2@     �G@     �B@     �N@      N@      &@      &@     �@@     �H@      @      (@     �C@      3@      7@     �A@     �A@     �S@      @       @      7@     �F@      @      @      8@      &@      .@      4@      :@     �H@      @      @      $@      @              @      .@       @       @      .@      "@      >@              �?     @S@      c@      "@      ,@     �^@      =@      q@      H@     �p@      W@      @      �?     @R@     �b@      @      ,@     �\@      5@      q@     �C@     pp@     �V@      @      �?     �B@      P@              @     �K@      ,@     �]@      8@      U@      D@       @              B@     @U@      @      @      N@      @      c@      .@     `f@     �I@       @              @      @      @              @       @       @      "@       @      �?                              �?      @              @               @      @       @                              @       @                       @       @              @              �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJw?�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @2=���J@�	           ��@       	                    �?�D_F-�@�           �@                          �;@�n�1v'	@W           ��@                           �?\C�KY�@�           �@������������������������       �pX+��v@�            ps@������������������������       ���h�@9           �~@                           �?�%���	@\             b@������������������������       ���v��@             F@������������������������       ����%�@?            @Y@
                          �4@�u�A��@�           @�@                            �?(�w���@w           Ў@������������������������       ��}0�&�?�            Ps@������������������������       ���*��@�           (�@                           �?ԯ;�+@*           ��@������������������������       �U>�7@�             r@������������������������       ������@�           ��@                           @���%+@�           �@                           �?����	@           ��@                           �?m��T�@�             m@������������������������       ��P��&@{             h@������������������������       ��ޏi��?            �C@                           �?��yw��	@s           ��@������������������������       ��~��~
@*           �}@������������������������       �F64�E@I            �]@                           �?�����@�            �p@                           �?�R*%�?6            �V@������������������������       �(����?"             I@������������������������       ��~{e���?            �D@                           @���@i            @f@������������������������       ���U�@             D@������������������������       �捽ZB&@S            @a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     �@      8@     @P@     �y@     �S@     ��@     �i@     h�@      x@      B@      "@      i@     0y@      *@     �E@     �q@      L@      �@     �a@     ��@     0q@      7@       @     @Y@     �`@      @      ;@      a@      6@     �^@      V@     �c@     ``@      0@      @     @U@      \@      @      9@      _@      .@     �]@     �R@     �`@      X@      ,@             �@@     �I@              @     �E@      @     �G@      D@     �B@      D@      "@      @      J@     �N@      @      4@     @T@      "@     �Q@     �A@      X@      L@      @      @      0@      4@      @       @      *@      @      @      *@      8@     �A@       @              @      @                      @      �?      @      @      &@      @              @      (@      ,@      @       @      @      @      �?       @      *@      =@       @      �?      Y@     �p@      @      0@     �b@      A@     (�@     �K@     �{@      b@      @              >@     @`@      @      @     �J@      @     {@      (@     `o@     �N@                      @      B@                       @             �c@      @     @S@      8@                      :@     �W@      @      @     �F@      @     Pq@       @     �e@     �B@              �?     �Q@     �a@       @      $@      X@      =@     �j@     �E@      h@     �T@      @              (@      E@      �?              7@      @     �V@      @      S@      ?@              �?      M@     �X@      �?      $@     @R@      7@     @^@     �B@      ]@      J@      @      (@     @U@     @e@      &@      6@      `@      6@     `n@      O@     �j@     �[@      *@      (@     �R@     �b@      $@      2@     �[@      5@     @`@      K@     `a@      W@      *@              0@     �D@      �?      @      8@              M@      1@      J@      4@                      0@      D@      �?      @      1@             �C@      0@      F@      1@                              �?                      @              3@      �?       @      @              (@      M@     �[@      "@      .@     �U@      5@      R@     �B@     �U@      R@      *@      (@      I@     �R@      "@      (@     @R@      4@      I@      8@     �R@     �N@      *@               @     �A@              @      *@      �?      6@      *@      (@      &@                      &@      3@      �?      @      3@      �?     @\@       @     �R@      3@                      @       @              �?       @             �L@              9@                              �?       @              �?      �?              B@              "@                              @                              �?              5@              0@                              @      1@      �?      @      1@      �?      L@       @     �H@      3@                       @      @              �?      @              $@       @      @      @                      @      (@      �?       @      ,@      �?      G@             �E@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��Ji#@�	           ��@       	                    �?�3��=@U           2�@                           �?��iTE�@�           ��@                          �4@1g'Td#@�            `y@������������������������       �&E��@�            �t@������������������������       �)�N(s<@,             R@                          �2@{�Q�
@�            `v@������������������������       �R���@�             h@������������������������       ��<:�9 @Z            �d@
                           @�(�4@~           t�@                            @:&|Z[�@8           @�@������������������������       �T�D#��@{           ��@������������������������       �n�V�G,	@�             s@                           @`*���v@F           ��@������������������������       ��w �Д@�            @u@������������������������       �$�thJ�?r             h@                            @���@7           ��@                           @c����p@�           �@                            �?�����M	@�           0�@������������������������       ��Qʳ�	@�            �r@������������������������       �·Gh�@�            �u@                          �8@�/�pKa@>           `@������������������������       �G�&���@�             q@������������������������       ���F6� @�            �l@                           @�"v��A	@Y           ��@                           �?�|��!	@7            @������������������������       �S־�j	@�             j@������������������������       �k�yڽ�@�            r@                          �9@�3��q@"            �P@������������������������       �	����@            �D@������������������������       �ڵ�{*A@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     8�@      >@     �L@     �x@      T@     ��@     `j@     ��@     �v@      7@       @     �[@     Pu@      (@      7@     �i@      8@     ��@     �U@     �~@     �c@      @              D@     �Y@       @      @     �N@      @     �t@      2@     �d@      A@                      2@     �J@       @      @     �A@      @     �g@      ,@     �P@      4@                      (@     �B@              @     �@@      @     �c@      *@     �K@      3@                      @      0@       @               @      �?      ?@      �?      (@      �?                      6@      I@               @      :@             �a@      @     @X@      ,@                      @      7@               @      3@              X@      @      C@      @                      0@      ;@                      @             �G@      �?     �M@       @               @     �Q@     �m@      $@      2@      b@      2@     @y@      Q@     �t@     �^@      @       @     �M@      f@      @      .@     @Z@      2@     �h@      P@     `c@     @W@      @      �?     �D@     �_@      @      @      N@      $@     �a@     �F@      Y@      O@       @      @      2@      I@      @      $@     �F@       @      K@      3@     �K@      ?@      @              (@      O@      @      @     �C@             �i@      @     �e@      =@                       @      D@      @       @     �A@             �]@      @     @Z@      9@                      @      6@              �?      @              V@      �?     @Q@      @              *@      e@      q@      2@      A@      h@      L@     pq@     @_@     `t@     @j@      0@      @      ]@     �e@       @      2@     �`@     �C@     �f@     �T@     `m@      b@      "@      @     �R@      Y@      @      0@      T@      @@      R@     �N@     �X@      X@      @       @      C@     �E@      @      $@      B@      $@      E@      A@      D@      C@      @       @      B@     �L@       @      @      F@      6@      >@      ;@     �M@      M@      �?      @      E@     �R@      @       @     �J@      @     @[@      5@      a@     �H@       @      @      6@     �D@       @      �?      <@      @      S@      @      Q@      4@       @              4@      A@      �?      �?      9@      �?     �@@      2@      Q@      =@              @     �J@     �X@      $@      0@     �M@      1@     �X@     �E@     �V@     @P@      @      @      G@     �T@      @      0@      J@      ,@     �S@     �C@     @V@      P@      @      @      5@      B@      @      &@      6@      @      @@      $@      ?@      @@      @              9@      G@      @      @      >@      $@     �G@      =@      M@      @@      @      @      @      1@      @              @      @      3@      @       @      �?                      @      0@                      @              (@      @       @                      @      @      �?      @              @      @      @      �?              �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Q�lhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Bb�f(@�	           ��@       	                   �;@g#���@           ��@                           �?\���t�@v           ĕ@                           �?��ė��@           0z@������������������������       ��Ý��X@�            `i@������������������������       �̡��7�@�             k@                          �4@�p���@g           p�@������������������������       ��K'�#U@           �z@������������������������       �m�0�@b           (�@
                           @�]��~	@�            �p@                          �<@p�+�@�            `m@������������������������       �S�R�F	@%             O@������������������������       ���d�7�@p            �e@                            �?�_8P|�@            �@@������������������������       �������@             4@������������������������       �H�j	"@             *@                          �4@;Q�x�@�           ��@                            �?�G�Q�@�           (�@                           @&/���@�           0�@������������������������       ��y�Ǩ@�            �r@������������������������       �o���@�            �w@                           @$��� @)           @~@������������������������       ���$|�@E             `@������������������������       ����p̎ @�            0v@                           �?+�� �m@�           �@                          �5@'t�J�@B            �@������������������������       �h�K��@A            �[@������������������������       �&ԕb@            y@                            �?8%�s�@i           �@������������������������       � ~���@�            0s@������������������������       ����9�s@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     `p@     Ȃ@      6@      I@     @}@     @T@     0�@     �j@     ��@     w@      @@      3@     @c@     �p@      &@      8@     �p@      J@     �m@     ``@     �n@      l@      :@      "@      _@     �l@      $@      4@     �m@      A@     �k@     �[@     �j@     �c@      6@             �F@     �Q@      @       @     �L@      @     �W@      9@     �S@     �@@      @              6@      8@      @      �?      @@      @     �J@      2@      <@      1@      �?              7@     �G@              �?      9@              E@      @     �I@      0@      @      "@     �S@     �c@      @      2@     �f@      ?@     �_@     @U@      a@     @_@      1@      @      >@      H@              @     �Q@      .@     @R@     �B@     �P@     �Q@      @      @     �H@     �[@      @      *@      \@      0@      K@      H@     @Q@     �K@      &@      $@      >@      C@      �?      @      >@      2@      0@      5@      =@     �P@      @      @      =@      ?@      �?      @      :@      0@      .@      (@      ;@     �O@      @      @      $@      @      �?              @      @      @              "@      (@      @      �?      3@      :@              @      5@      $@      $@      (@      2@     �I@      �?      @      �?      @                      @       @      �?      "@       @      @               @              �?                      �?       @              "@       @      @              �?      �?      @                      @              �?                      �?               @      [@     �t@      &@      :@     �h@      =@     ��@     �T@     �@      b@      @             �H@     �e@       @      ,@     �Q@       @     �~@      @@     �p@      O@                      A@     �[@      �?      @     �D@             @o@      0@      g@      C@                      ;@     �K@                      2@             @X@      &@     �Q@      3@                      @     �K@      �?      @      7@              c@      @     @\@      3@                      .@     �O@      �?      $@      >@       @      n@      0@     �T@      8@                      �?      0@      �?      @      0@             �H@      $@      3@      (@                      ,@     �G@              @      ,@       @      h@      @     �O@      (@               @     �M@      d@      "@      (@      `@      ;@     0s@     �I@     �n@     �T@      @       @      ?@     @S@      �?      "@     �O@      "@      _@      6@      ^@     �H@      @              �?      2@                      "@      @      C@              >@      @       @       @      >@     �M@      �?      "@      K@       @     �U@      6@     �V@      F@      @              <@     �T@       @      @     @P@      2@     �f@      =@     �_@     �@@      �?              (@      K@       @      �?      ;@      (@     �U@      2@      R@      6@                      0@      =@      @       @      C@      @      X@      &@     �K@      &@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJX6�DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�t��Sl@�	           ��@       	                    �?��RO_�@V           4�@                           �?�`��G@�           ��@                            @h���1�@�            �x@������������������������       ����"��@�            �r@������������������������       ���ŏc@>            �W@                            @����Z�@�            u@������������������������       ��v��{�@�            �m@������������������������       ���r�g@<             Y@
                          �1@��A@�           �@                          �0@i�	��^@�             w@������������������������       �f��Τ@E             \@������������������������       �ЏĦ~�@�             p@                           @1S
bگ@�           $�@������������������������       ��N���@�           @�@������������������������       ���G)/@�            x@                          �8@�o�ΰ�@H           ��@                           �?SP
�@�           ��@                           @��l�\@�             v@������������������������       ��\�g@�            s@������������������������       �
�&�7@            �H@                            @Y�t�E�@           �z@������������������������       �f�6��@�            �s@������������������������       ��ᜍ�@J            �\@                           �?#S���?	@U           ��@                          �9@���0
@C           �~@������������������������       �4��@7             V@������������������������       ��}j�
@           `y@                           @v^�Y�@           {@������������������������       �ӑǭ�@�            pw@������������������������       �#�c��@%             M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �p@     P�@      <@      O@     @|@     @W@     ��@      o@     �@     �u@      >@      $@     @Z@     �t@      (@      7@     �k@      G@     Є@     �\@     �@     �c@       @              @@     �X@              @      J@       @     �r@      8@     �f@      A@       @              1@      I@              @     �A@       @     �d@      0@      U@      2@       @              @      E@              �?      @@      @     @`@      ,@      P@       @       @              *@       @               @      @       @     �A@       @      4@      $@                      .@     �H@              �?      1@             �`@       @     @X@      0@                      .@      A@                      $@              W@      @      R@       @                              .@              �?      @              E@       @      9@       @              $@     @R@      m@      (@      3@      e@      C@     �v@     �V@     �t@     �^@      @       @      ,@      H@              @      B@      �?      `@      4@      V@      =@                      @      2@                      "@             �I@              0@      (@               @       @      >@              @      ;@      �?     �S@      4@      R@      1@               @     �M@      g@      (@      0@     �`@     �B@     �m@     �Q@      n@     @W@      @       @     �H@      `@      @      ,@     �X@     �@@     @Y@     �P@     �_@      S@      @              $@      L@      @       @     �@@      @      a@      @     �\@      1@      �?      @     @d@     �o@      0@     �C@      m@     �G@     �s@     �`@     Pr@     �g@      6@              T@     �`@      @      2@     �\@      5@     �d@      8@     �a@     �R@      "@             �@@     �L@      �?       @     �D@              X@      @     �P@      B@      "@              @@     �F@              @     �A@             �U@      @      K@     �@@      "@              �?      (@      �?      @      @              "@              (@      @                     �G@     @S@       @      $@     @R@      5@     �Q@      1@     �R@      C@                      D@      I@       @      "@     �F@      .@     �N@      ,@     �N@      2@                      @      ;@              �?      <@      @      "@      @      ,@      4@              @     �T@      ^@      *@      5@     �]@      :@     �b@     �[@      c@     @]@      *@      @     �H@      Q@      (@      *@     �R@      .@      K@     �R@      G@     @Q@      (@               @      (@      @              2@      �?      @      :@       @      @      @      @     �D@      L@      "@      *@     �L@      ,@     �H@      H@      C@     �P@       @             �@@      J@      �?       @     �E@      &@     �W@      B@     �Z@      H@      �?              2@     �F@               @     �C@      "@      V@      <@     �W@      F@      �?              .@      @      �?              @       @      @       @      &@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJYȾ:hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @F0�(M@�	           ��@       	                    �?��b��@�           �@                           �?>�3�@,           �@                           �?����>@�            Pr@������������������������       ���N�@T             a@������������������������       �0-�ȓ�@i            �c@                           @k��6E�@o           ��@������������������������       �~���� @           �x@������������������������       �e2kHm�@h            �b@
                          �4@O�K�+�@�           Ğ@                          �1@�v��@           �@������������������������       ���\��@�            @p@������������������������       �x*�:@o           ��@                          �<@j�ː=�@�           <�@������������������������       ���*ȶ�@U           Ѝ@������������������������       ��$W���@_            �b@                           @���@�           T�@                          �?@�����@           H�@                           �?C��Ǥ�@           8�@������������������������       �+8���@t             f@������������������������       ��f�l�@�           ��@                           @�0N��@             A@������������������������       �U�}�6@             6@������������������������       ��[���@             (@                           @����n@�            �p@                           �?���*�O @S            �`@������������������������       ���+Z{F�?;            @X@������������������������       ��k��X@            �B@                           �?�ai �@W            �`@������������������������       ��.[��� @*             P@������������������������       �4v�2�@-            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     ps@     �@      =@      I@     �{@     �Q@     ��@     @k@     ��@     `x@      >@      $@     �k@     �w@      (@      ?@     �s@      L@     ��@      a@     ��@     �p@      9@      @     �M@     �]@       @       @      U@      @     �q@      3@     �g@      M@      @      @     �A@     �G@      �?      �?     �I@      @     �D@      *@      N@      B@       @      @      1@      3@                      5@              ;@      @      >@      0@                      2@      <@      �?      �?      >@      @      ,@      $@      >@      4@       @              8@     �Q@      �?      �?     �@@      @     �n@      @     @`@      6@      @              5@     �E@                      3@      @     �g@      @     @Y@      *@      @              @      <@      �?      �?      ,@      �?     �L@      @      =@      "@       @      @      d@     `p@      $@      =@     �l@     �H@     @}@     @]@     �y@     `j@      2@             �H@     �Z@      @      @      U@      @     �q@      >@     @i@     �U@      @               @     �A@              �?      (@       @     �\@      @     �O@      3@                     �D@     �Q@      @      @      R@      @     �e@      9@     `a@     �P@      @      @      \@     �c@      @      6@      b@     �E@     �f@     �U@     �i@     @_@      ,@      @      U@     �a@      @      5@     �]@     �A@     �e@     �Q@     �g@     �W@      $@              <@      *@              �?      :@       @      @      0@      .@      ?@      @      ,@     �V@     �d@      1@      3@     �`@      ,@     Pp@     �T@     `g@     @^@      @      ,@     �T@     �a@      *@      .@     �\@      *@     �b@     @S@     �Z@     @[@      @      $@     �R@     @a@      *@      &@      [@      *@     �b@      S@      Z@      Z@      @       @      *@      ?@      �?      @      5@             �E@      @      >@      8@      �?       @      O@     �Z@      (@      @     �U@      *@     �Z@     �Q@     �R@      T@      @      @      @      @              @      @                      �?      @      @              @      @      �?               @      @                      �?       @      @                      @      @               @                                      �?       @                      "@      8@      @      @      2@      �?     �[@      @      T@      (@                      @      (@               @       @             �Q@      @      =@      �?                      �?      @              �?      @             �M@       @      6@      �?                      @      @              �?      @              (@      @      @                              @      (@      @       @      $@      �?      D@             �I@      &@                              �?      @               @      �?      1@              =@      @                      @      &@      �?       @       @              7@              6@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @ӀǹS\@�	           ��@       	                    �?o����@�           ��@                           �?2v��%@�           ��@                          �;@�G��U@�             t@������������������������       ��'q�r@�            �p@������������������������       � bbh]�@             I@                           �?M�\8�@�            �u@������������������������       �Tɽh@�            @p@������������������������       ��`\��@?            �V@
                          �5@�Ʌ\Q	@�           ��@                          �0@�X�)}@�           ��@������������������������       ����&O@!            �I@������������������������       �j:(�@�           ��@                           �?�]�~�	@           ��@������������������������       �i�5�a�	@2            �T@������������������������       �O:�`i	@�           X�@                           �?d͗B@           �@                          �4@w�W0d@e           @�@                          �0@���?�             t@������������������������       �vz��V�?%            �I@������������������������       ��n��U��?�            �p@                          �7@�p��2�@�            �l@������������������������       ���b*�@F             _@������������������������       ��XE�;@E            �Z@                           @0����T@�           L�@                           �?�%k�ֲ@p            �f@������������������������       �oR�ܯ@'            @P@������������������������       ��0���@I            @]@                           @�
� �@H           �@������������������������       �M��^��@�           ��@������������������������       �q:�+@�            pp@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     0t@     �@      <@     �J@     �{@     �R@     ��@     �l@     ��@     �w@      :@      2@     �l@     u@      6@      D@     �q@      K@     �w@      h@     �x@     0q@      9@             �P@     �V@       @      &@      T@      @     `g@      9@      b@     �K@      @              ;@      D@       @      @     �C@      @     @X@      .@     �M@      >@                      7@      @@       @      @     �@@      �?     �W@      &@     �J@      2@                      @       @               @      @      @      @      @      @      (@                      D@      I@              @     �D@             �V@      $@     �U@      9@      @              @@     �E@              @     �A@              N@       @     �K@      3@       @               @      @                      @              >@       @      ?@      @      �?      2@      d@     �n@      4@      =@     �i@      H@     `h@      e@     @o@     �k@      6@      &@     �P@      ]@      @      $@     @X@      2@     �\@      P@     �b@      X@      @               @      4@              �?      @               @      @      @      @              &@     @P@      X@      @      "@      W@      2@     �Z@     �N@     �a@     �V@      @      @     �W@     ``@      ,@      3@      [@      >@      T@      Z@     @Y@      _@      2@      @      $@       @              @      $@      @       @      *@      .@      "@       @       @      U@     �^@      ,@      *@     �X@      ;@     �S@     �V@     �U@     �\@      0@      �?     �W@     �m@      @      *@     `c@      4@     ��@      C@     �x@     �Z@      �?              :@     �R@              �?      ?@      @     @p@      $@     �_@      4@                      4@      ;@              �?      "@              f@      @     @R@      &@                              "@                       @              ;@              &@       @                      4@      2@              �?      @             �b@      @      O@      "@                      @     �G@                      6@      @      U@      @     �J@      "@                       @     �C@                      .@       @     �C@              6@      @                      @       @                      @       @     �F@      @      ?@      @              �?     @Q@     @d@      @      (@      _@      0@     �t@      <@     �p@     �U@      �?      �?      "@     �@@              "@      4@      @      K@      "@      >@      &@              �?      @      ,@               @      &@      @      "@      @      $@      @                       @      3@              @      "@      @     �F@      @      4@      @                      N@      `@      @      @      Z@      $@     �q@      3@     �m@      S@      �?             �F@     �W@       @      �?      O@      @     �l@      *@     `e@     �B@      �?              .@     �A@      @       @      E@      @      I@      @     �P@     �C@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�٦`hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @���@�	           ��@       	                    �?��i�%p@q           j�@                          �<@�*�O@�           �@                           �?0aj��a@w           ��@������������������������       ����@           �z@������������������������       ����V7.@h             f@                          @@@�\\Fq�@3            �W@������������������������       ��+7d@*            �S@������������������������       � �rN@	             0@
                           �?��	�	@�           ��@                           �?�a��Mf	@�           (�@������������������������       �[�o7��@            z@������������������������       �� xڲ�	@�           P�@                            @�;��{N@           �z@������������������������       �����B%@�             r@������������������������       ���.��@R            �a@                          �4@x�uc��@I           P�@                            �?�%��@S           0�@                          �1@.����?�            �i@������������������������       ���q��V�?5            �T@������������������������       ��iΉ @W            @^@                           @��d
T�@�           Ѕ@������������������������       ��dLg@E           P@������������������������       ���"��@�            �h@                            @���h��@�           p�@                          �7@8 $��@�           (�@������������������������       �}x�8|�@�            �s@������������������������       ��WQ @�            �t@                           @�؄F�@U             a@������������������������       ���xh1s�?*            �R@������������������������       ���-��@+             O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �s@     ��@      A@     �H@     �|@     �S@     t�@     `g@     �@     �v@      7@      $@      m@     �s@      <@      ?@     `t@      P@     �y@     �b@     �x@      o@      2@              S@     �W@      @      "@      S@      @      g@      @@     �c@      N@      @              Q@     @T@      @      @     �P@      @     �f@      7@     �a@      ?@       @              L@     �P@      @      @     �J@       @      \@      6@     �U@      5@       @              (@      ,@                      ,@      @      Q@      �?     �K@      $@                       @      *@              @      "@              @      "@      .@      =@      �?               @      (@              �?      @              @      "@      $@      =@      �?                      �?              @      @               @              @                      $@     �c@     �k@      8@      6@     @o@     �M@     �l@     �]@     `m@     �g@      .@      $@     �_@     �b@      8@      0@     �f@      F@     �a@      T@     �d@      b@      .@              :@     �M@      @      @     �R@      (@     �T@      =@      N@      O@      @      $@      Y@      W@      5@      *@     �Z@      @@     �M@     �I@      Z@     �T@      $@              >@     @Q@              @     @Q@      .@      V@      C@     �Q@      F@                      3@      D@              @      M@      "@      K@      >@     �J@      6@                      &@      =@              �?      &@      @      A@       @      2@      6@               @     @U@     �k@      @      2@      a@      .@     ��@     �B@     �y@     �[@      @              E@     �[@      @      "@     �H@       @     �y@      .@     @j@     �I@                      @      3@              �?      (@             �]@      @     �A@      $@                              @              �?      @              L@      �?      *@      @                      @      0@                       @             �O@      @      6@      @                      C@     �V@      @       @     �B@       @     @r@      &@     �e@     �D@                      5@      O@      �?      @      3@       @     �l@      @     @`@      =@                      1@      =@       @      @      2@              P@      @     �F@      (@               @     �E@     �[@      @      "@      V@      *@     `l@      6@      i@      N@      @       @      D@     �X@      �?      @     �R@      *@     �e@      1@      d@      J@      @              *@     �O@      �?      @      @@       @     �Y@      @     @P@      2@      @       @      ;@      B@              @     �E@      @     @R@      *@      X@      A@                      @      &@       @       @      *@              J@      @     �C@       @       @              �?       @                      @              C@              7@       @       @               @      "@       @       @      @              ,@      @      0@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���&hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ؼ��?@�	           ��@       	                    �?�
�Ȼ@�           ��@                            @QߔՒ/@4           `~@                           �?��A�W0@�            �q@������������������������       ���'�^@O             `@������������������������       ���=]�@g            `c@                          �=@
0�-�%@~            @i@������������������������       �J��K�@t             g@������������������������       �H �D�J@
             1@
                           @�+��,@�           Ѕ@                          �=@)i�|@�            �p@������������������������       ���ܿO@�             p@������������������������       ��ڇ8�E@             (@                           @�B�J?Z @           �z@������������������������       ���_:e�?�            `l@������������������������       �r�̜*�@�             i@                           @l%�+�	@�           R�@                          �9@����	@�           �@                           �?��D���@�           ��@������������������������       �1�$��@           x�@������������������������       �K���`�@�            �v@                           �?�y��7�	@�            0x@������������������������       ��@� :�@             A@������������������������       ���:�j	@�            v@                          �1@��[o�@�           ��@                          �0@�	ҍ�E�?~            `i@������������������������       ��\K�%��?!             I@������������������������       �&l$���?]             c@                           @�;l�@F           �@������������������������       �ea�עk@�            @j@������������������������       �k~�;@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     ��@      A@     �K@     �}@     �S@     �@     `l@     ��@     �u@      6@       @     @T@     `d@      @      ,@      Z@      @      z@      H@     q@     �P@      @       @     �I@     @T@      @      (@     �L@       @     �Y@      <@     @Z@     �D@       @       @      6@      H@      @              @@       @     �M@      &@     @S@      :@       @       @       @      8@      @              ,@       @      =@      "@      6@      0@                      ,@      8@                      2@              >@       @     �K@      $@       @              =@     �@@              (@      9@             �E@      1@      <@      .@                      <@      ?@              @      6@              E@      0@      <@      &@                      �?       @              @      @              �?      �?              @                      >@     �T@               @     �G@      @     �s@      4@      e@      :@       @              5@     �C@                      3@      @     @X@      &@     @P@      *@      �?              3@     �C@                      1@      @      X@      @      P@      *@                       @                               @              �?      @      �?              �?              "@     �E@               @      <@      �?     `k@      "@     �Y@      *@      �?              @      5@                      @      �?     `b@              E@      @                      @      6@               @      5@              R@      "@     �N@      "@      �?      1@     @k@     �w@      ?@     �D@     pw@     �Q@     �@     `f@     �@     `q@      2@      0@     �a@     �n@      3@      ;@     �p@      O@      n@      c@     �j@     `h@      .@       @     @Z@     �h@      .@      6@     �i@      9@     �i@     �Y@     @f@     �`@      $@       @     �U@      a@      ,@      .@     `e@      1@     @\@     �R@     �Z@     �W@      $@              2@     �O@      �?      @      B@       @     �V@      =@     �Q@     �B@               @      B@     �F@      @      @      N@     �B@     �B@      I@     �B@     �O@      @      @      @      @              �?      @                      @       @      @      @      @     �@@      C@      @      @      L@     �B@     �B@     �E@     �A@     �M@       @      �?     @S@     �`@      (@      ,@      [@      "@      w@      :@     �r@     �T@      @               @      9@               @      &@             �V@       @     �P@      @                      �?      @                                      8@              2@      @                      �?      6@               @      &@             �P@       @      H@                      �?     �R@     �[@      (@      (@     @X@      "@     Pq@      8@      m@     �S@      @      �?      =@      @@       @              9@      @     �J@      @     �E@      ,@       @              G@     �S@      $@      (@      R@      @      l@      5@     �g@     @P@      �?�t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�A�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �? FjV4B@�	           ��@       	                    �?���*�O	@            <�@                           �?Q �^��@:           �~@                          �2@�7f���@o            �e@������������������������       �i�t�7@            �H@������������������������       �0x�R��@U             _@                          �6@�)�m�@�            �s@������������������������       ���9m��@t            �f@������������������������       ���*�@W             a@
                           @��_&��	@�           ��@                           �?L����p	@�            @l@������������������������       �ĎmZ��@=            �V@������������������������       �6�T$x%	@T            �`@                          �>@QAz9�	@5           �@������������������������       �t2�D��	@            �@������������������������       �A5�ԂQ@'            �O@                           �?��j��@�           ��@                          �=@��0�&�@�           @�@                           @�݅ʇU@�           ��@������������������������       �;Y�� @V           ��@������������������������       �`5�U@|            �g@������������������������       ��;�\�Z@             3@                           @$ �g�@�           H�@                          �5@��7��@�           x�@������������������������       ��4���@�            @x@������������������������       �/����@�            �r@                          �<@6�w"�@'           �@������������������������       �,1)G�@           ��@������������������������       ��!h�R�@            �B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     �s@     ؁@      @@     �N@     �z@     �R@     8�@     �k@     H�@     �u@      ;@      1@     �f@     �n@      5@      C@      l@      H@      p@     �`@     �l@      i@      5@             �I@     �R@       @      "@     �H@      @     �[@      @@     @X@     �N@      �?              .@      :@                      .@              H@      @      E@      5@                              @                      @              5@      @      (@       @                      .@      3@                      &@              ;@      @      >@      3@                      B@     �H@       @      "@      A@      @      O@      :@     �K@      D@      �?              :@      5@      �?       @      ,@      @      I@      (@      =@      7@                      $@      <@      �?      @      4@              (@      ,@      :@      1@      �?      1@     @`@     �e@      3@      =@      f@     �F@     @b@      Y@     ``@     �a@      4@      @      <@      6@      �?      @     �C@      $@      ,@      =@      C@      >@      @       @       @      $@              �?      7@      @      &@       @      2@      &@       @      @      :@      (@      �?       @      0@      @      @      5@      4@      3@      @      &@     �Y@     �b@      2@      :@      a@     �A@     �`@     �Q@     @W@     �[@      ,@      $@     @V@     `a@      1@      :@      a@      ?@     �_@     @P@     �U@     @X@      *@      �?      *@      &@      �?                      @      @      @      @      *@      �?              a@     @t@      &@      7@     �i@      ;@     p�@     @V@     (�@      b@      @              >@     �V@       @      �?     �I@      @     �t@      (@     �g@      =@       @              >@     @V@       @      �?      G@      @     �t@      @     @g@      ;@      �?              =@      N@                      =@      @      o@      �?     �a@      3@                      �?      =@       @      �?      1@             �T@      @      F@       @      �?                      �?                      @                      @      @       @      �?             �Z@     @m@      "@      6@     `c@      6@      |@     @S@     pv@     �\@      @              G@     �`@       @      (@     �M@      0@     �e@      I@      `@     �P@       @              *@     �U@       @      @      >@       @      ^@      9@     �Q@      ;@       @             �@@     �G@               @      =@       @     �J@      9@     �L@     �C@                     �N@     @Y@      @      $@      X@      @     Pq@      ;@     �l@     �H@       @              J@     �X@      @      "@     �T@      @      q@      ;@     `l@     �G@       @              "@       @       @      �?      ,@              @              @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�zZj@�	           ��@       	                   �8@�����~	@�           �@                           �?��F��@�           ��@                            @C+u(({@�            `x@������������������������       �b/KX{�@�            `h@������������������������       ��C��|v@w            `h@                           �?�K�>w:@�           ��@������������������������       ��
}n�r@�            0p@������������������������       ��S�7v@           �z@
                            @�
"^�}
@=           �@                            �?:,�	s�	@�            �r@������������������������       ���JL�
@�            �p@������������������������       ��+*��q@            �C@                          �9@6<���{
@�            @j@������������������������       �+#:��@             E@������������������������       ��Z@��
@k             e@                           �?��h�@�            �@                           �?�I�k�F@�           h�@                           @�=`D+�@�            �x@������������������������       ��5�@�@c             b@������������������������       ���x L�@�            �o@                            �?Xh�8�@�            �s@������������������������       �	5��� @<            �Y@������������������������       �X����� @�             k@                          �4@�H�@�           �@                          �1@k�Ս�@�           @�@������������������������       �ww���f @�            �o@������������������������       �S��e@�@P           X�@                           @�e�f�Q@�           ؈@������������������������       �*��Ǥ2@�            �j@������������������������       ��%:Z�@u           8�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     Pr@     ��@      >@      M@     �{@     �U@     �@     �l@     �@     w@      <@      5@     �e@     `o@      8@      D@     �k@      H@      l@      a@     @n@     @h@      5@      @     �^@     �d@      *@      7@     �c@      8@     �g@      S@     �f@     @\@      @       @     �A@     �S@       @      "@      O@      @     �Q@      ;@     �C@     �H@      @              4@     �F@               @      <@      @      ?@      6@      2@      7@      @       @      .@      A@       @      @      A@      @     �C@      @      5@      :@      �?      @     �U@      V@      @      ,@      X@      2@     �]@     �H@     �a@      P@      @              =@      @@      �?      @      =@      @      N@      1@     �I@      <@      �?      @      M@      L@      @      $@     �P@      &@     �M@      @@      W@      B@       @      .@      I@      U@      &@      1@      O@      8@     �A@      N@      N@     @T@      ,@      @      <@      F@       @      @     �D@      6@      5@      A@     �B@     �J@      @      @      7@      D@       @      @      <@      3@      3@      A@      @@     �G@      @      �?      @      @                      *@      @       @              @      @               @      6@      D@      "@      $@      5@       @      ,@      :@      7@      <@      @              @      1@      @       @      @                      @      @               @       @      2@      7@      @       @      2@       @      ,@      4@      2@      <@      @             @^@     ps@      @      2@     `l@      C@     �@     @W@     x�@     �e@      @              <@     @T@      �?      @     �I@      &@     �s@      "@     �f@     �A@      �?              *@      I@              @      A@      @     �f@      @     @S@      ;@                      @      5@                      $@      @     �J@      @      =@      2@                      @      =@              @      8@      @     �_@      @      H@      "@                      .@      ?@      �?              1@      @     �`@       @      Z@       @      �?                      3@      �?              @       @     �E@      �?      =@      �?      �?              .@      (@                      (@      @      W@      �?     �R@      @                     @W@     �l@      @      ,@      f@      ;@      |@      U@     �w@     �a@      @              <@     �Y@      �?      @      N@      @      s@      B@      h@      R@                       @      =@              �?      $@             �_@      &@      N@      ,@                      :@     @R@      �?      @      I@      @     �f@      9@     �`@      M@                     @P@      `@      @       @      ]@      7@      b@      H@      g@      Q@      @              7@      D@              @      @@      (@      6@      8@     �B@      1@       @              E@      V@      @      @      U@      &@     �^@      8@     �b@     �I@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��kFhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����)@�	           ��@       	                    �?ԟ�.Q@           ��@                          �;@��S�@*            @                            �?���@           �z@������������������������       ���Yt�@R            �_@������������������������       �`�{J�5@�            �r@                            �?�+��@(            �P@������������������������       �Qӯmi�@             E@������������������������       ��[�z�A@             9@
                          �5@w�em��@�           ؇@                           @I?�YL @E           p�@������������������������       ���󄍇�?�            �x@������������������������       ��᯲�o@V            �_@                          �=@����6@�            �m@������������������������       �rIv)@�            �i@������������������������       �����X@             >@                           @:��{#@�           ��@                           �?�xxt	@�           (�@                          �8@��p�@�             y@������������������������       ��E�$B`@�            �r@������������������������       ��?�9�@?            �X@                           �?e�\�F�	@�           ��@������������������������       ��㱇e
@�           ��@������������������������       ���c3�@           z@                          �4@DG�"��@�           P�@                           @�u��@Y           (�@������������������������       ��g��@�            �u@������������������������       ���GZt@l             e@                           �?�h^�N@q           x�@������������������������       �Xk��J@�            pq@������������������������       �������@�            �s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     ��@      9@      L@     �{@      U@     <�@     �g@     ��@     0v@     �@@      @      Q@      f@      @      "@     @[@      "@     P}@     �D@     0q@     �W@       @      @     �C@      T@       @      @     �N@      @      _@      8@     �V@     �N@      �?              @@     �P@       @      @      K@      �?      ]@      6@      U@     �F@      �?               @      2@              �?      0@              ?@      @     �A@      *@      �?              8@     �H@       @      @      C@      �?     @U@      2@     �H@      @@              @      @      *@              �?      @      @       @       @      @      0@              @      @      @                      @      @      �?       @      @      0@                      @      @              �?      @              @              @                              =@     @X@      �?      @      H@      @     �u@      1@      g@     �@@      �?              1@     @Q@              @      =@             �p@      &@     @]@      $@      �?              0@      H@              �?      5@             �j@      @     @V@      @                      �?      5@               @       @              K@      @      <@      @      �?              (@      <@      �?              3@      @      S@      @     �P@      7@                      $@      ;@      �?              *@      @     @R@      @      O@      ,@                       @      �?                      @      �?      @      @      @      "@              0@     �n@     �v@      6@     �G@     �t@     �R@     Ё@     `b@     �@     Pp@      ?@      .@     �e@     �l@      1@     �B@     �l@     �O@     @j@     �]@     �o@     �e@      ;@              8@      L@       @      &@     �R@       @      O@      <@     �S@     �J@      @              3@      G@       @      &@      J@      @      J@      1@      P@     �A@                      @      $@                      6@      @      $@      &@      .@      2@      @      .@     �b@     �e@      .@      :@     @c@     �K@     �b@     �V@      f@     �]@      6@      .@      Z@     �W@      ,@      1@     �W@     �F@      R@     �L@     �[@     �T@      4@             �F@      T@      �?      "@      N@      $@      S@     �@@     @P@      B@       @      �?     �R@     �`@      @      $@     �Y@      (@     �v@      =@     �q@     @V@      @              ?@      P@      �?      @      ?@      @     @j@      "@     �`@     �@@                      9@      H@      �?      �?      ;@      �?     �`@      @     �U@      9@                      @      0@               @      @       @     �S@      @      G@       @              �?     �E@     �Q@      @      @      R@      "@     �b@      4@     @c@      L@      @      �?      3@     �A@              @      A@      @      O@      @     �S@      =@      @              8@      B@      @              C@      @      V@      ,@     �R@      ;@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJÛ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?(��T�[@�	           ��@       	                   �4@�v�Z@'           H�@                           @MF��@�           ��@                           �?[,�7�@�            0t@������������������������       ������l@T            �`@������������������������       ����@x            �g@                           @���:�?�            0u@������������������������       ��纳��?�            `o@������������������������       ����	�@>             V@
                           �?\ �cP@w           ��@                            �?���y9@�             s@������������������������       �+���|�@o             e@������������������������       �zB3�@Q             a@                          �=@� �"��@�            �p@������������������������       ��`N��@�            `n@������������������������       �J����@             7@                           @"ϚGL@�           �@                           @�C�nL @�           L�@                            @`�f�Wt	@K           ��@������������������������       ���fcr@�            `v@������������������������       ��̯�
@o            �e@                            �?���f`@g           L�@������������������������       �������@           �z@������������������������       ��(Lچ@M           ��@                           !@K9*�k	@�            u@                           @��+	@�            �s@������������������������       �ypZi�	@~            �g@������������������������       ��A��Kl@K            @^@������������������������       ���c�{@             9@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        7@     s@     �@      =@     �M@     �~@     @V@     X�@     @k@     Ј@      u@      7@             @X@      f@       @      (@     �]@      @     0|@      E@     �p@     �N@      @             �A@     @T@              @     �J@      �?     �r@      .@      c@      9@                      5@      E@              �?      D@      �?      [@      &@      U@      .@                      @      .@                      8@      �?     �E@      "@      =@      @                      ,@      ;@              �?      0@             @P@       @     �K@       @                      ,@     �C@              @      *@             �g@      @      Q@      $@                       @      =@                      @             @b@      �?     �K@      @                      @      $@              @       @              E@      @      *@      @                      O@     �W@       @       @     @P@      @     `c@      ;@     @\@      B@      @             �G@      K@      �?       @      E@             �I@      1@     �K@      <@      @              :@      :@      �?      @      :@              2@       @      B@      3@      @              5@      <@               @      0@             �@@      "@      3@      "@                      .@     �D@      �?              7@      @      Z@      $@      M@       @                      .@      D@      �?              4@      @     @X@      @     �K@      @                              �?                      @      �?      @      @      @       @              7@      j@     �v@      ;@     �G@     Pw@     �T@     @�@      f@     ��@     Pq@      4@      0@      g@     �s@      8@      F@     pt@     �Q@     p@     �`@      ~@      m@      &@      (@     �D@     �N@      @      (@     �V@      ;@     @T@     �D@     @Y@      J@      @      @      :@     �B@              "@     �O@      .@      M@      ;@     �R@      D@      @      @      .@      8@      @      @      ;@      (@      7@      ,@      :@      (@      @      @     �a@     �o@      2@      @@     �m@      F@     `z@      W@     �w@     �f@      @       @      >@     �L@              @     �O@       @     @_@      :@     @R@      D@               @     @\@     �h@      2@      9@     �e@      B@     �r@     �P@      s@     �a@      @      @      8@     �H@      @      @      G@      &@     �H@     �E@     �H@      F@      "@      @      4@     �H@      @      @     �D@      @     �H@     �E@      F@     �C@      "@      @      *@     �@@               @      <@      @      7@     �@@      2@      7@      @              @      0@      @      �?      *@              :@      $@      :@      0@      @              @                              @      @                      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�:>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@��=��>@�	           ��@       	                    �?Pͥ��(@b           ��@                            @�5��@�           8�@                           @�$̏�@(           �~@������������������������       ��־�@l            @g@������������������������       ��h/����?�             s@                           �?4�M���@n            `g@������������������������       ��]��I�@7            �V@������������������������       �R���?7            @X@
                           @���	��@�           �@                          �1@���T�i@z           ��@������������������������       ��Xa:�@p            �f@������������������������       ��pg��
	@
           �y@                           @.}"���@R           P�@������������������������       �؀���V@�            0q@������������������������       ����:�@�            pq@                          �;@���bm@*           N�@                           @��T�@           ��@                           �?��D�r�@g            �@������������������������       �a��)P	@�            pv@������������������������       �%c���[@w           �@                           @p�5@m@�           @�@������������������������       ���OK�@�           P�@������������������������       ��8�@(             O@                          �?@"/�"j	@           �{@                          �=@MP�]8�@�             u@������������������������       ����@�            @i@������������������������       �\��
@@S            �`@                            �?W�Jk��	@A            �Z@������������������������       �"B��[�@             G@������������������������       �æ�Vp@#            �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     0r@      �@      ;@      O@     p|@     �T@     (�@     �k@     H�@      u@      ?@       @      X@     �m@      "@      8@     @d@      2@     ��@     �U@     0w@      b@      "@             �A@      S@              @      H@      @     `s@      ,@     �c@      @@      �?              7@      M@               @     �A@             �k@      &@      ^@      3@      �?              &@      4@              �?      :@             �L@       @      K@       @      �?              (@      C@              �?      "@             �d@      @     �P@      &@                      (@      2@               @      *@      @     �U@      @      B@      *@                       @      *@               @      @      @      >@      @      *@      (@                      @      @                      @             �L@              7@      �?               @     �N@      d@      "@      4@     �\@      .@     `v@      R@     �j@     @\@       @       @     �C@     �U@      @      ,@     @V@      (@     �_@     �O@     �S@      Q@       @              "@      @@       @       @      6@             �I@      1@      @@      ,@               @      >@     �K@      @      (@     �P@      (@      S@      G@     �G@      K@       @              6@     @R@      @      @      9@      @     �l@      "@      a@     �F@                      (@     �E@      �?              1@      @     �[@      @      L@      :@                      $@      >@      @      @       @             @^@       @      T@      3@              *@     `h@     �u@      2@      C@     Pr@     @P@     �v@      a@     `y@     �g@      6@      @     @c@     q@      *@      9@     �l@      E@     @t@      Z@     Pt@     @`@      3@      @     �]@     @e@      "@      4@     �c@      A@      `@     @V@      c@     �Q@      &@       @      A@      M@      @      @     �K@      *@      Q@      :@     �J@      >@      @      @      U@      \@       @      ,@     �Y@      5@      N@     �O@      Y@      D@      @              B@     �Y@      @      @     @R@       @     �h@      .@     �e@      N@       @             �A@      W@      �?      @     @P@      @     @f@      (@      e@      L@      �?              �?      &@      @               @      @      2@      @      @      @      @       @     �D@     �Q@      @      *@     �O@      7@      E@      @@     @T@     �N@      @      @      8@      N@      �?      *@      H@      2@     �A@      4@     @P@      G@      �?      @      0@      @@      �?      @      4@      "@      3@      $@      K@      >@                       @      <@              @      <@      "@      0@      $@      &@      0@      �?      @      1@      &@      @              .@      @      @      (@      0@      .@       @              "@      @                      @      @      �?      @      @      "@       @      @       @      @      @              "@              @      @      *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�u�~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?,Pso�)@�	           ��@       	                   �8@�[�@           ��@                           �?L4V(�@�            �@                           �?�\L��+@�            �w@������������������������       �L��B4@h            `f@������������������������       �1�����@~            �i@                           �?�d��`@�           �@������������������������       �,z��� @�            x@������������������������       � 1K.g@�             p@
                            �?%�"\7-@�            @m@                            �?����u@M            @\@������������������������       �[q\3�,@)             J@������������������������       ���@$            �N@                          �>@�{evQ�@L            @^@������������������������       �PpO��@@             Y@������������������������       �w�Sڲ�@             5@                           @.��Z@�           ��@                          �9@���h5	@�           ��@                           �?\��)Sq@�           `�@������������������������       �D���:�@           ��@������������������������       ������@�            �u@                            �?YY
@�             v@������������������������       ���^���	@>             Y@������������������������       ��I�<�	@�            �o@                           @ �/e5@�           ��@                           @��̙�L@�            �@������������������������       ��0���@�           X�@������������������������       ��q�|F�@             9@                            �?�?�%��@�            0t@������������������������       �F�$��@7            �U@������������������������       �3�2�@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     �@      ?@      L@     �|@     �Q@     ��@     @j@     ��@      v@      >@       @     @U@     �d@      @      &@      \@      .@     0|@      ;@     Pr@     �U@      @             @Q@      ^@      @      @      U@      @     �y@      5@     @n@      K@      @             �E@      H@       @      @      C@      @      X@      (@     �X@     �@@      @              5@      7@       @       @      9@      @     �G@      @      @@      .@      @              6@      9@              �?      *@             �H@      @     �P@      2@       @              :@      R@       @      @      G@      @     �s@      "@     �a@      5@      �?              1@     �G@              @      A@      @      i@      @      Q@       @                      "@      9@       @              (@             @\@      @     �R@      *@      �?       @      0@      F@              @      <@       @     �D@      @     �I@     �@@      �?       @      @      7@              @      "@      @      $@      @      5@      <@      �?       @       @      (@                       @      @      @       @      (@      "@      �?              @      &@              @      @       @      @      �?      "@      3@                      $@      5@              �?      3@      �?      ?@      @      >@      @                      $@      3@              �?      ,@      �?      <@      @      8@                                       @                      @              @              @      @              ,@     �l@     �u@      ;@     �F@     �u@     �K@     x�@     �f@     X�@     �p@      7@      ,@     �d@      j@      4@      ?@      l@      F@     �j@     �b@     �p@     �d@      5@      @     @_@      g@      &@      <@     @f@      3@     @g@     @Z@     @k@     �Z@      $@      @     �Y@     �]@      "@      9@      `@      .@     �[@     �Q@     �c@      T@      $@              6@     �P@       @      @      I@      @      S@     �A@     �N@      :@               @     �D@      9@      "@      @     �G@      9@      :@      F@     �J@      N@      &@       @      @      @      @      �?      3@      @      $@      3@      .@      &@      @      @     �B@      5@      @       @      <@      3@      0@      9@      C@     �H@      @              P@     �a@      @      ,@      _@      &@     �u@      A@     �q@     �X@       @             �F@     @Y@      @      @     �T@      @     pq@      :@     @i@     �J@       @             �D@     @Y@      �?      @     �S@      @     @q@      6@      i@     �H@       @              @               @              @       @      @      @      �?      @                      3@      D@      @      &@     �D@      @      Q@       @     �T@      G@                      @      @              �?      "@              ;@      @      1@      0@                      (@     �A@      @      $@      @@      @     �D@      @     @P@      >@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJݢ�MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @xr��t�@�	           ��@       	                   �6@�R �3@           8�@                          �1@�:Z	��@~           <�@                            �?�uu��@-           �~@������������������������       �R�)r�@�            `v@������������������������       �*���T�@Q             a@                           @�q1Y@Q           ��@������������������������       �6��1c@�           H�@������������������������       ��:M[T@�           ��@
                           �?�wO�6�@�           4�@                            �?n��ua@�            �r@������������������������       ����D�d@B            �Z@������������������������       �fίF��@r            `h@                          �:@��%��%	@�           ��@������������������������       ����	�	@           |@������������������������       ��Fx��@�            �q@                           �?�騾�-@�           ��@                          �=@,�7��(	@�           0�@                          �5@�'p���@�           x�@������������������������       �?#`�ּ@�            �r@������������������������       ��<.�.5	@�            Pr@                          �>@1�)���@%            �K@������������������������       �b!	;<L@             1@������������������������       �x�{��@             C@                           @�ρ+��@           pz@                          �3@�$�f�N@f            �c@������������������������       ���B��@(             N@������������������������       �>��)�G@>            @X@                           @ۊc��@�            �p@������������������������       �f={�d@P            ``@������������������������       ��JA�`�@Z            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     `s@     0�@      =@     @P@     �}@     @W@     p�@      n@     P�@     �v@      ;@      @     �j@     �w@      2@      C@     Pt@     �Q@     h�@      e@     P�@     �p@      6@      @      ^@      n@      &@      4@     �e@      8@     p�@      W@     0x@     �`@      $@      @      5@      H@               @     �I@       @      j@      3@     �X@      B@      @      @      0@     �D@               @     �@@       @     @b@      *@     �P@     �A@                      @      @                      2@              O@      @      @@      �?      @      �?     �X@      h@      &@      2@      _@      6@     �w@     @R@      r@     �X@      @      �?     �N@     �T@      @      1@     @U@      0@     �\@      L@      ]@     �M@       @              C@     �[@      @      �?     �C@      @     �p@      1@     �e@     �C@       @       @     �W@     �a@      @      2@     �b@     �G@     �c@     @S@     �h@     ``@      (@              :@      H@      �?              ;@      "@     �M@      $@     �S@      D@      @              $@      4@      �?              ,@      @      .@      @      @@      @       @              0@      <@                      *@      @      F@      @     �G@      A@      �?       @     @Q@      W@      @      2@     �^@      C@      Y@     �P@      ^@     �V@      "@              D@     �N@      @      ,@      P@      6@     �Q@      G@     �S@     �D@       @       @      =@      ?@      @      @     �M@      0@      =@      5@     �D@      I@      �?       @     �W@     @e@      &@      ;@     `b@      6@      l@     �Q@      h@      X@      @       @     @T@     @Z@       @      3@     @Z@      3@     �S@      G@     �Y@     @Q@      @      @     @R@     �W@      @      *@     @W@      3@     @S@     �F@     �Y@     �M@      @      @      =@      E@      @      @     �J@      @     �I@      ,@     �N@      @@      �?              F@     �J@      @      $@      D@      *@      :@      ?@     �D@      ;@      @      @       @      $@      �?      @      (@              �?      �?      �?      $@                      @                      @      @              �?                      @              @      @      $@      �?      �?      @                      �?      �?      @                      ,@     @P@      @       @      E@      @     `b@      9@     @V@      ;@                      @      <@       @      @      2@      �?      H@      2@      4@      (@                      �?      "@              @      �?              8@       @      "@      @                      @      3@       @              1@      �?      8@      $@      &@      "@                      "@     �B@      �?      @      8@       @     �X@      @     @Q@      .@                      @      1@               @      "@      �?      M@      @      ?@      �?                      @      4@      �?      �?      .@      �?     �D@              C@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJom4hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�N��]@�	           ��@       	                   �4@"Tr�I@�           ��@                           @��"��@C           @�@                          �2@�a��ģ@�            �@������������������������       �
Ͼ��@�            �w@������������������������       ������@�            pt@                            �?�C��&9@v           ��@������������������������       ��
�x�@�            �w@������������������������       ��g&Eh��?�            �j@
                           �?�`�C�@�           �@                          �8@gp��9�@	           `z@������������������������       ��j$@�             o@������������������������       �e酃@k            �e@                          �<@8#�>A6	@�           ��@������������������������       ��r5c��@N           ��@������������������������       �G�ǜa@W             a@                           @zy�ɿ�@�           ȑ@                           �?�?��@#            �@                           �?g�\×�@�           h�@������������������������       �._H]M@            �h@������������������������       ����cO�	@0           �~@                          �3@=O�JB@t            �f@������������������������       �ʌ���/@*            �P@������������������������       ��V�b�@J            @]@                           �?��)m�$@�            �p@                           �?��]" @E             [@������������������������       ��Dn�� @&             O@������������������������       ���E���?             G@                          �7@ƕZ�9�@p            @d@������������������������       �:�:w��@O             ]@������������������������       �,҄���@!             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     pq@     ��@      <@     �N@     �}@     �U@     ��@     `k@     Ј@     pv@      A@      @     �f@      y@      1@     �F@     �t@     �P@     �@     `b@     ��@      p@      5@             �Q@     @d@      @      @     @^@      &@     @|@      G@     �r@     �]@      @              N@      V@      @      @     �V@      &@      h@     �C@     �`@     �R@      @              =@      H@                      E@      @     �`@      1@     @P@      A@      @              ?@      D@      @      @      H@      @      M@      6@     �Q@     �D@       @              $@     �R@       @       @      ?@             0p@      @     `d@     �E@      �?              @     �C@       @       @      9@             �b@       @      ]@      B@                      @     �A@                      @             @[@      @     �G@      @      �?      @     �[@     �m@      (@      C@      j@      L@     �q@     @Y@     �p@     @a@      .@              ;@     @Q@      �?      @      F@      "@      _@      4@      X@      9@       @              4@      B@      �?      @      =@      �?     �V@      @     �J@      @                      @     �@@                      .@       @     �@@      *@     �E@      3@       @      @      U@      e@      &@     �@@     �d@     �G@      d@     @T@     �e@     @\@      *@      @     �Q@     @c@      &@      >@     �a@      =@     �b@     �Q@     �d@     @T@      (@      �?      ,@      .@              @      6@      2@      (@      &@       @      @@      �?       @     �X@     �e@      &@      0@     �a@      4@     �o@      R@     @l@     �Y@      *@       @     @V@     �b@      $@      *@     @]@      2@     �a@      Q@     @d@     �T@      (@       @     �Q@     �\@      $@      $@     �Y@      .@     @W@      J@     �_@      R@      (@              5@     �D@              �?      5@             �H@      "@      E@      *@               @     �H@     �R@      $@      "@     @T@      .@      F@     �E@      U@     �M@      (@              3@      A@              @      .@      @     �G@      0@      B@      $@                      @      "@              @       @              ;@      @      .@       @                      0@      9@                      *@      @      4@      &@      5@       @                      "@      :@      �?      @      :@       @     @\@      @      P@      5@      �?              �?      "@              �?      @       @     �N@      @      5@      @                      �?      @              �?      @              ?@      �?      .@      @                              @                       @       @      >@      @      @                               @      1@      �?       @      5@              J@             �E@      1@      �?              @      *@      �?              (@              F@              >@      $@      �?              @      @               @      "@               @              *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��{8hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @GXd�m@�	           ��@       	                    �?��:l	@�           �@                           �?��z-�@-           x�@                            �?���� c@.           @}@������������������������       �m�.i�6@�            pu@������������������������       ����� ��?M            @_@                          �6@V^E�l�@�            �y@������������������������       �u<-@�            0q@������������������������       ��\	�@X             a@
                          �:@�q���@�           $�@                           @뺌[�@           ��@������������������������       ���ΤD	@           ��@������������������������       ��U�U@           8�@                          �=@�C6 ��@�            `r@������������������������       �+�M:e�@s            �e@������������������������       ���k��@D            �]@                           �?2�b�A@�           D�@                           �?��SO]t	@�           �@                          �8@D�Y�5�@j            �c@������������������������       �*	#�@T            @^@������������������������       �db.@             B@                           �?����0�	@L            �@������������������������       ��8AM�	@{            �e@������������������������       �*���T	@�            Pu@                           @���J�@            {@                          �1@��\M��@j             d@������������������������       ��ǒ?���?             8@������������������������       ��/0&^@Z             a@                          �3@�íL�@�             q@������������������������       ��ε%�<�?E             ^@������������������������       �~�*�0@d             c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     h�@      >@      N@     @{@     �U@     Ȏ@     �k@     p�@     0w@      =@      &@      i@     �x@      3@      F@     `r@      O@     H�@     @b@     (�@     p@      2@      �?      D@     �`@       @      @     �P@      @     t@      :@      l@     �H@      @      �?      0@     �P@      �?      @     �A@      @      h@      3@     �Y@      9@              �?      .@      E@      �?      @      =@      @      `@      .@     @T@      8@                      �?      9@                      @       @      P@      @      6@      �?                      8@     @P@      �?       @      @@      �?      `@      @     �^@      8@      @              1@     �F@                      $@             �Y@      �?      V@      (@                      @      4@      �?       @      6@      �?      :@      @      A@      (@      @      $@      d@     �p@      1@     �C@     `l@      L@     �z@      ^@     @x@      j@      *@      @     �`@     �l@      ,@      C@     �e@     �@@     y@     �W@     �u@     �c@      (@      @     �V@     @`@      @      ;@     �\@      =@     �`@     @R@      \@     @X@      $@              E@     �X@       @      &@     �M@      @     �p@      5@     @m@     �N@       @      @      =@      C@      @      �?      K@      7@      7@      :@      E@      I@      �?      @      .@      7@       @             �@@      "@      ,@      $@      >@     �A@                      ,@      .@      �?      �?      5@      ,@      "@      0@      (@      .@      �?      &@     �Y@     �c@      &@      0@     �a@      8@      n@     �R@      i@     �\@      &@      &@     @T@      X@       @      $@     @X@      7@     �V@     �L@     �Y@     �U@      &@              0@      ;@               @      1@       @      D@      1@      7@      *@                      &@      6@              �?      &@       @     �C@       @      3@       @                      @      @              �?      @              �?      "@      @      @              &@     @P@     @Q@       @       @      T@      5@      I@      D@     �S@     �R@      &@      @      8@      =@      @      @      9@      "@      $@       @      2@      A@      @      @     �D@      D@      @      @     �K@      (@      D@      @@     �N@      D@       @              5@     �O@      @      @     �F@      �?     �b@      1@     �X@      ;@                      "@      A@      �?       @      2@              F@      .@      7@      ,@                      �?      "@                                      "@              @                               @      9@      �?       @      2@             �A@      .@      2@      ,@                      (@      =@       @      @      ;@      �?     �Z@       @      S@      *@                      @      $@                      @              N@             �B@      @                      "@      3@       @      @      4@      �?      G@       @     �C@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ3�yRhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���
^@�	           ��@       	                   �1@�<���@[           ��@                           �?fd+�I@�           ��@                           �?f"�V4E@m             e@������������������������       �RwXSSw@5            @R@������������������������       ���i�'@8            �W@                           �?g�޻V@           p{@������������������������       ����<�@�            �l@������������������������       ���:t��?�             j@
                           �?L���e�@�           ė@                           @�c�j=�@M           ��@������������������������       ����@�            �p@������������������������       ���c��?�            `p@                           @޵�한@�           �@������������������������       �qDk��B@6           @�@������������������������       ����S�@N            @^@                           �?�{f�@M           �@                          �8@[��ӱ�	@%           H�@                          �6@�/���@�             x@������������������������       ��:�r@X            `a@������������������������       �Ҵ��[@�            �n@                           �?6_M:�u	@>           8�@������������������������       ��Az�۟@c             e@������������������������       ��#/up	@�            �u@                           �?9�X�@(           ��@                            �?���aa@�            �k@������������������������       �s> +�O@             E@������������������������       �R����g@q            `f@                           @�g�!�j@�           ��@������������������������       ��U�I&@x            �e@������������������������       ��Z�@$           @~@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pr@     p�@      A@     �Q@     �|@     @S@     ��@     �j@     @�@     �w@      4@      @     �Z@     �s@      *@      >@     �k@      >@     ��@     �U@     �@     �d@      $@      �?      <@     @T@      �?      @      J@       @     �n@      &@     @a@     �C@       @      �?      (@      ?@      �?      �?      ;@       @      =@      @     �C@      5@              �?       @      *@      �?              (@       @      .@       @      *@      (@                      $@      2@              �?      .@              ,@       @      :@      "@                      0@      I@              @      9@             @k@      @     �X@      2@       @              (@      :@              @      2@             �\@      @      D@      $@                      @      8@                      @              Z@      �?     �M@       @       @      @     �S@     `m@      (@      9@      e@      <@     �x@     �R@     �v@     �_@       @              @@     �Q@       @       @      >@      @     �h@      1@      a@      B@      �?              9@      <@       @       @      8@      @     �N@      ,@     �S@      <@      �?              @      E@                      @       @      a@      @      M@       @              @     �G@     �d@      $@      7@     @a@      7@     `h@      M@     �l@     �V@      @      @      D@      b@      $@      3@      ^@      2@     `e@     �J@      k@     �R@      @       @      @      5@              @      2@      @      8@      @      .@      0@      @      &@     @g@     @n@      5@      D@     �m@     �G@     �s@      `@     �t@     �j@      $@      "@     @X@     �a@      *@      @@     �`@      @@      X@      U@     @`@      `@       @       @     �J@     �O@      @      0@      L@      *@     �J@      3@     �P@     �B@      @       @      <@      @@       @      @      &@      @      ,@      "@      ,@      1@                      9@      ?@      @      (@     �F@      @     �C@      $@      J@      4@      @      @      F@      T@       @      0@     @S@      3@     �E@     @P@      P@     �V@      @       @      *@      7@       @       @      7@      @      8@      *@      =@      ?@       @      @      ?@     �L@      @      ,@      K@      .@      3@      J@     �A@      N@      @       @     @V@     �X@       @       @     �Y@      .@      k@     �F@     �i@     �U@       @              "@      :@      �?              $@      @     @T@      $@     �P@      *@      �?                      @      �?              �?              2@      �?      (@       @      �?              "@      4@                      "@      @     �O@      "@      K@      &@               @      T@     @R@      @       @     @W@      &@      a@     �A@     `a@     �R@      �?              <@      7@              @      >@      @      9@      .@      8@      3@      �?       @      J@      I@      @      @     �O@      @     �[@      4@     �\@     �K@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Z[$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?VY�8�@�	           ��@       	                    �?4�>D��@           �@                           �?���3�@           �{@                          �5@t��@f            �d@������������������������       � \�Rz@9            �W@������������������������       ���KUL�@-            �Q@                            �?z!J��=@�            pq@������������������������       �����@,             O@������������������������       �O��#r�@�             k@
                            @M�4'@�           X�@                          �4@�=::��@�           `�@������������������������       ��ӗ˃��?�            �v@������������������������       �;���@�            p@                           �?x�%Q;��?[            �c@������������������������       ���xю�?4            �U@������������������������       ��ӫv/d�?'             R@                           �?u ��k�@�           �@                          �9@S���	@�           �@                           �?����>	@�           x�@������������������������       ��:��&k@�            �r@������������������������       �c���	@8           0~@                           �?	�,���	@�            �r@������������������������       �������@2            �T@������������������������       �J����"
@�            `k@                           @�͛ߟ@�           �@                          �3@��JX�@           �z@������������������������       ��8�~��@c            `b@������������������������       �����[@�            pq@                            �?���@�           p�@������������������������       �M�x�_�@�            0p@������������������������       �Ρ�O`�@:           Ȍ@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     `r@     ��@      =@      H@     p|@     �L@     @�@     `l@     (�@      u@      ;@       @     �V@     �`@      @      *@     �[@      @      ~@     �E@     Pq@     �O@       @       @     �I@      M@      �?      @     @Q@      �?      X@      >@     @V@     �C@      �?       @      5@      2@                      0@              K@      @      C@      $@      �?              @      "@                      @              C@      @      >@      @               @      1@      "@                      &@              0@      �?       @      @      �?              >@      D@      �?      @     �J@      �?      E@      9@     �I@      =@                      "@      ,@                      (@              $@       @      *@       @                      5@      :@      �?      @     �D@      �?      @@      7@      C@      ;@                     �C@     @S@       @      @      E@      @      x@      *@     �g@      8@      �?              C@     �R@       @      @      >@      @      r@      (@     �a@      7@      �?              4@     �@@              @      &@             �i@      @     @R@      &@      �?              2@     �D@       @              3@      @     �U@      @     @Q@      (@                      �?      @              �?      (@             �W@      �?      G@      �?                      �?      �?              �?       @              K@              5@      �?                               @                      @              D@      �?      9@                      5@     �i@     Py@      :@     �A@     �u@     �J@     ��@      g@     ��@     q@      9@      5@      ^@     �c@      .@      3@     @f@     �B@     @]@     �Z@     @b@     �b@      3@      0@     �U@     �]@      "@      ,@     �a@      .@      X@      P@     �]@     @V@      .@              5@      K@      @      @     �I@      �?     �J@      5@     �G@     �D@       @      0@     @P@      P@      @      "@     �V@      ,@     �E@     �E@      R@      H@      *@      @      A@     �C@      @      @      B@      6@      5@      E@      ;@      N@      @              @      "@       @              *@      @       @      *@       @      7@              @      ?@      >@      @      @      7@      3@      *@      =@      3@     �B@      @              U@      o@      &@      0@     �d@      0@     �{@     �S@     �y@      _@      @              6@     @W@      @      @     �I@      @      U@     �G@     �U@      =@       @              @      <@                      "@             �I@      ,@      ?@       @                      0@     @P@      @      @      E@      @     �@@     �@@     �K@      5@       @              O@     `c@       @      *@     �\@      $@     pv@      ?@     �t@     �W@      @              2@     �@@      @              4@       @     �T@      &@      P@      9@                      F@     �^@      @      *@     �W@       @     @q@      4@     �p@     �Q@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJU�b<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@�h@�	           ��@       	                   �1@�y(�$,@0           ��@                           �?g��|�@r           0�@                           �?�ٍn�v@o            �d@������������������������       ��"��,@6             U@������������������������       ��N��k�@9            �T@                           @!' ��@           �y@������������������������       �8�0�5�@�            @t@������������������������       ���ESc��?9            �V@
                           @��h�@�           �@                           �?�վ~�T@�           ��@������������������������       �F���@�            u@������������������������       �)�N��	@           p�@                          �4@-&�R�\@�            �@������������������������       �즟���@9           �}@������������������������       ��e�S��@�            �l@                           �?m��@�            �@                           �?i�4<@�             y@                          �;@��R�`�@�            �h@������������������������       �*���4�@V            �`@������������������������       �߸����@*             P@                          �9@W"�K��@y            �i@������������������������       ���x��@@            �Z@������������������������       ���K�[@9            �X@                           @m�i�2	@�           p�@                           �?[o%�	@�           ��@������������������������       ��z�=�
@R           �@������������������������       �f]c��@\            @b@                           @9�:��@�            �u@������������������������       �a5�.{�@�            �k@������������������������       ��o}��s@N            @_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@      �@     �B@     �K@     }@     �U@     x�@     �j@     @�@     Pw@      :@       @     �d@     pv@      ,@      A@     Pp@      B@     ��@     @[@      �@     �i@      (@              @@     �T@      �?      @     �F@      @     �m@      2@     �]@      D@                      (@      <@      �?      �?      9@      @      D@      @      =@      5@                      @       @                      *@      @      @@       @      .@      @                       @      4@      �?      �?      (@               @      @      ,@      ,@                      4@      K@              @      4@             �h@      &@     @V@      3@                      4@     �D@               @      4@             `b@      @     @R@      0@                              *@               @                     �I@      @      0@      @               @     �`@     Pq@      *@      =@      k@     �@@     �@     �V@     �z@     �d@      (@       @     @[@      i@      "@      8@     �c@      ?@     �m@     �T@     �k@     @^@      (@              <@      I@              @      ;@       @     @X@      (@      V@      <@      �?       @     @T@     �b@      "@      4@     �`@      =@     �a@     �Q@     �`@     @W@      &@              8@      S@      @      @     �L@       @     `q@       @      j@     �F@                      0@     �E@      @      @      ;@             �h@       @     �a@      A@                       @     �@@      �?      �?      >@       @     �S@             �P@      &@              @     �b@      g@      7@      5@     �i@     �I@     �k@      Z@     @p@     �d@      ,@      �?      A@     �K@      @      $@      I@      @     @V@      .@     �X@     �A@       @      �?      ;@     �@@       @      $@     �A@      @      4@      *@      <@      7@       @              .@      8@       @      @      <@              2@      &@      5@       @       @      �?      (@      "@              @      @      @       @       @      @      .@                      @      6@      @              .@      @     @Q@       @     �Q@      (@                      @      &@      @              @             �D@              =@      @                              &@                       @      @      <@       @      E@      @              @      ]@     @`@      1@      &@     @c@     �F@     �`@     @V@      d@     �`@      (@      @     �S@     �U@      ,@      "@     �X@     �D@      P@     �R@     �T@     �W@      &@      @      P@     �P@      ,@      "@     �R@      =@     �G@      O@      P@     �P@      $@              .@      4@                      7@      (@      1@      *@      2@      ;@      �?      �?     �B@     �E@      @       @      L@      @     @Q@      ,@     �S@      C@      �?      �?      :@      9@                      C@      @      L@      @     �I@      0@      �?              &@      2@      @       @      2@      �?      *@      "@      <@      6@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�0+x8@�	           ��@       	                     �?{D��o"@           ��@                           �?AWq�y@�           8�@                          �<@���k�@�            Px@������������������������       ����Y,R@�            �v@������������������������       �t�����?             6@                          �8@v!rt�@�             t@������������������������       ���F�@�            p@������������������������       ��?� N@*            @P@
                          �2@�M<�@b           @�@                           �?=6��O�@~            `h@������������������������       �r�Ơ@>            �V@������������������������       ���Ô�@@             Z@                          �=@���g��@�            Pv@������������������������       ��Hx��S@�            �t@������������������������       ���9��@             8@                           @�?�h�;@�           ��@                          �2@����@�           $�@                           @mR%�@l           ��@������������������������       ��g��&@�            �w@������������������������       ��ꃛf�@r            �f@                            �?�?I�x~@K           ��@������������������������       ���թ��@,           �~@������������������������       �&�S@           ē@                          �4@s�Y�4�	@�            �t@                          �0@A�}c�@H            @Z@������������������������       �l ����?             &@������������������������       �)�]UWy@A            �W@                           @�gU���	@�            �k@������������������������       ��*E ��@`            `c@������������������������       �ݶ���@.             Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �p@      �@      4@     �P@     @|@     �V@     �@      j@     �@     �v@     �@@             �S@      g@              0@     �W@      $@     �|@      C@     �r@     �T@       @              F@      Z@               @      I@      @     �n@      8@     @e@      N@       @              3@      M@              @      E@      @     �a@      (@     @R@      B@                      3@      J@              @      E@       @      a@      (@      R@      :@                              @                              �?      @              �?      $@                      9@      G@               @       @       @      Z@      (@     @X@      8@       @              0@     �C@                      @             �X@       @     @S@      ,@                      "@      @               @      @       @      @      @      4@      $@       @             �A@     @T@               @      F@      @     �j@      ,@     �_@      7@                      &@      "@              @      ,@             @X@      @      E@      (@                      @      @                      @              F@      @      6@      @                       @      @              @       @             �J@      @      4@      @                      8@      R@              @      >@      @     �]@      @     @U@      &@                      8@      Q@              �?      5@      @     �\@      @     �T@      &@                              @              @      "@              @              @                      1@      g@     px@      4@     �I@     `v@      T@     ��@     @e@     @@     pq@      ?@       @     @c@     `u@      1@      I@     @s@      N@      �@     �a@     �|@     �n@      6@              :@     �Q@       @      @     �K@              h@      D@     �^@      H@      �?              (@      I@       @      @      G@             �_@      3@     @X@      ;@                      ,@      5@              �?      "@             �P@      5@      :@      5@      �?       @      `@     �p@      .@      G@     �o@      N@      t@      Y@     @u@     �h@      5@      @     �B@     @R@              .@     �Q@      1@     @Z@      E@     @R@      J@      @      @     �V@     �h@      .@      ?@     �f@     �E@     �j@      M@     �p@     @b@      .@      "@      ?@     �H@      @      �?      I@      4@      L@      >@     �B@     �@@      "@      �?      @      $@              �?      .@      �?      =@      @      4@      ,@      @                                              �?              "@      �?                              �?      @      $@              �?      ,@      �?      4@      @      4@      ,@      @       @      ;@     �C@      @             �A@      3@      ;@      9@      1@      3@      @       @      1@     �@@      �?              6@      2@      (@      5@      @      .@      �?              $@      @       @              *@      �?      .@      @      $@      @      @�t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJe�g,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?y)�".@�	           ��@       	                     �?s���OI	@�           0�@                          �:@�����n@,           p}@                          �5@e�S�7�@�            w@������������������������       �@b޹<y@�            �h@������������������������       �(NΙ�@g            `e@                           �??����w	@>            �Y@������������������������       ���Z@             <@������������������������       ��)=�E	@+            �R@
                          �?@E+p�e�	@�           ԑ@                           �?\ܨ�D	@�           А@������������������������       �� uD6@�            �t@������������������������       ���i#w�	@�           H�@                            @���O@"            @P@������������������������       ��f���0@             3@������������������������       �4r�V��@             G@                          �3@�q"��@�           ��@                          �1@%���@o           `�@                           @���\� @           �{@������������������������       ��W�&� @�            @v@������������������������       �4z-��� @?            �U@                           @�<��x@Q           ��@������������������������       �(M��@�            0u@������������������������       �fX�C4@�            �g@                          �=@���+�;@=           Ĕ@                           @�C�/��@           D�@������������������������       �s����@R           ؀@������������������������       ����X�@�           ��@                           @�CU�*	@8             X@������������������������       �O���	@&            @P@������������������������       ��:X��@             ?@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      q@     �@      B@     �L@     �}@     �R@     L�@     �j@     x�@     �t@      ;@      7@     �c@     �l@      7@     �A@     �p@     �D@     @o@     @`@     0p@     �e@      :@      �?      B@      P@      @      $@     @U@      &@     �R@      H@     @U@      G@      @              @@      L@       @      @     �P@       @     �N@     �C@     �Q@      =@      @              1@     �@@              �?      :@      �?     �C@      ,@      G@      3@       @              .@      7@       @      @      D@      �?      6@      9@      9@      $@      @      �?      @       @       @      @      3@      "@      ,@      "@      ,@      1@      �?      �?      �?      @                       @       @      @       @      @                              @      @       @      @      &@      @      "@      @       @      1@      �?      6@      ^@     �d@      3@      9@     �f@      >@     �e@     �T@     �e@     �_@      4@      1@     �Y@     �d@      1@      3@     `e@      ;@     �e@     @S@     �d@     �]@      4@              >@      F@      @      @      I@      �?     @T@      6@      O@      ;@      @      1@     @R@     @^@      *@      *@     @^@      :@     �W@     �K@      Z@      W@      0@      @      1@      �?       @      @      $@      @              @       @       @                       @                       @      �?      @                      @       @              @      "@      �?       @      @      "@                      @      @      @              �?      ]@     �s@      *@      6@      j@      A@     Ȉ@     �T@     `�@     �c@      �?              B@     �_@      �?      @      P@              z@      4@      o@     �J@                      .@      J@              @      ?@             `m@      "@      S@      5@                      ,@     �D@              �?      >@             `g@      @      P@      .@                      �?      &@              @      �?              H@      @      (@      @                      5@     �R@      �?      @     �@@             �f@      &@     �e@      @@                      &@      K@      �?      @      3@              ^@      @     �\@      *@                      $@      4@                      ,@             �N@      @     �M@      3@              �?      T@     �g@      (@      .@      b@      A@     �w@      O@     0s@     �Z@      �?      �?      R@     �f@      &@      &@     @`@      >@     �v@      I@     @r@     �V@              �?     �D@     @W@              @      Q@      4@     @_@      ?@     @]@     �B@                      ?@      V@      &@      @      O@      $@     �m@      3@     �e@      K@                       @      "@      �?      @      ,@      @      *@      (@      .@      .@      �?               @       @      �?      @      $@      @      "@      &@      @      &@      �?              @      �?                      @              @      �?      &@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?"�4�k@�	           ��@       	                    �?C�/@i�@           ��@                          �<@�{�U<@>           �@                            �?l�5�?@           �|@������������������������       �/���@�            @o@������������������������       ���&�x@�             j@                           �?���%�@&            �K@������������������������       ��1�ZP�@             8@������������������������       �c�/F@             ?@
                          �=@�2�A?�@�           (�@                           �? S7f|@�           x�@������������������������       �/�.��-@            y@������������������������       ���<4� @�            �s@������������������������       ����^ @             6@                            @�F���R@�           Ƥ@                           @<��)�@�           ��@                           @CS׮�@�           ܜ@������������������������       ��,��gF	@Q           ��@������������������������       ��KkZ%�@H            �@                           �?�V���@             �G@������������������������       ���}�@
             .@������������������������       ��+Dk�@             @@                           �?��%�@�           �@                           �??�Ya�@�            @s@������������������������       ��J}DR/	@x             g@������������������������       ��E�"@S            �^@                          �4@Q�&�@-           �|@������������������������       ��u(ۻ�@u            �e@������������������������       ���%�`@�            �q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        9@      s@     Ё@      ;@      G@     �|@      T@     p�@     �m@     x�@     �w@      <@      �?     @V@      f@       @      "@     �\@      "@     �{@      F@     pq@     �T@      @      �?     �G@      W@       @       @     @R@      @     @Y@      >@      Y@     �I@      @      �?      D@     @T@       @       @      P@      @     �X@      8@      X@     �A@      @      �?      5@     �B@       @      @      @@              J@      ,@      P@      2@      @              3@      F@              @      @@      @     �G@      $@      @@      1@                      @      &@                      "@               @      @      @      0@                      @       @                      @              �?               @      @                       @      @                      @              �?      @       @      (@                      E@     @U@              �?      E@      @     @u@      ,@     `f@      @@      �?              C@     @U@              �?     �C@      @     u@      @     `f@      >@      �?              7@      L@              �?      9@       @     �h@      @     @S@      ,@                      .@      =@                      ,@      �?     @a@      �?     �Y@      0@      �?              @                              @       @      @       @               @              8@      k@     �x@      9@     �B@     pu@     �Q@     ��@     `h@     �@     `r@      7@      (@      a@     �q@      ,@      ;@     `m@      H@     �y@      c@     �v@     �h@      ,@      &@      `@     �q@      ,@      ;@     �l@     �F@     @y@     �a@     `v@     @h@      $@      "@      U@     �a@      "@      1@      b@      C@      ]@     �[@      `@     @\@      $@       @      F@     `b@      @      $@     @U@      @      r@      =@     �l@     @T@              �?       @                              @      @      @      *@      @       @      @                                                       @       @      @      �?       @      �?      �?       @                              @      �?      @      @       @              @      (@     @T@     �Z@      &@      $@      [@      7@     �^@      E@     �a@     �X@      "@       @      ?@      G@      "@      @      ?@      "@      L@      &@      L@     �F@      @       @      =@      >@      @       @      ;@      @      .@      @      9@      >@      �?               @      0@      @      �?      @      @     �D@      @      ?@      .@       @      @      I@      N@       @      @     @S@      ,@     �P@      ?@     �U@     �J@      @      @      $@      2@              @      :@      @     �D@      &@     �D@      ,@      @      �?      D@      E@       @      @     �I@      $@      9@      4@      G@     �C@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�OshG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��I)�V@�	           ��@       	                     �?���y@           ��@                          �8@-����@�            pu@                          �0@Y�^] �@�            0q@������������������������       ���mbl��?            �@@������������������������       ��� {�G@�            @n@                           �?Ĥ K2X@+             Q@������������������������       ��!:��@            �A@������������������������       ��5>�g@            �@@
                          �<@W�#��@*           ��@                          �4@Ƨnam�@�           Ȉ@������������������������       ���:�{�@           �{@������������������������       ��&a^�@�            �u@                            �?>ML@+            �O@������������������������       �L��A�@             <@������������������������       �l�B&��@            �A@                           @�a�U@�           4�@                          �3@����u~	@�           h�@                            @�F}�R@           p{@������������������������       �Fr@�            �p@������������������������       ���{�@k             e@                           @�15m��	@�           ��@������������������������       �9)�8��	@d           ��@������������������������       �ǧ��9�@U            �a@                           @I��Llw@�            �@                           @5hh�Q@�           ��@������������������������       �cY��@�            �@������������������������       ��3���@�            �s@                          �4@��Ιi@             =@������������������������       �=*,I�R @             &@������������������������       �u���#�?             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@      9@     �I@     0}@     �S@      �@     �j@     0�@     0u@     �E@       @     @R@     `e@      �?       @     �Y@      $@     �z@      @@     pr@      S@      �?       @      $@     �H@              @      5@      @     �^@      @     �X@      7@      �?              @      B@              @      3@      �?     �[@      @     �T@      ,@                       @      @                      @              1@               @      �?                      �?      =@              @      .@      �?     �W@      @     @T@      *@               @      @      *@                       @      @      (@       @      .@      "@      �?       @      @      @                      �?       @      @      �?       @      @                      @      "@                      �?      @      @      �?      @      @      �?             �O@     �^@      �?      @     �T@      @      s@      ;@     �h@     �J@                     �M@     @[@      �?       @     �R@      @     �r@      6@     �g@      C@                      1@     �K@               @     �E@       @     �g@      0@     @X@      7@                      E@      K@      �?              ?@       @      [@      @     �V@      .@                      @      *@              �?       @               @      @      "@      .@                      �?      @              �?                      @      @      @      (@                      @      $@                       @              @       @      @      @              0@      n@     px@      8@     �E@     �v@      Q@     Ȁ@     �f@     ��@     pp@      E@      0@      d@     @n@      7@      9@     `n@     �J@      i@      b@     �n@      e@      C@      @      :@     �S@       @      @      O@       @     �X@      8@     @S@      J@      @              1@     �H@       @             �E@       @      P@      4@     �F@      ;@       @      @      "@      =@              @      3@      @     �A@      @      @@      9@      �?      (@     �`@     �d@      5@      5@     �f@     �F@     �Y@      ^@     @e@     @]@     �A@      "@     @]@     �a@      3@      5@     �c@      E@     �W@     �V@     �c@     �Y@      :@      @      2@      6@       @              6@      @       @      =@      &@      ,@      "@             �S@     �b@      �?      2@     @^@      .@      u@     �C@     �r@     �W@      @              R@     `b@      �?      0@     @\@      .@     �t@     �B@     0r@     @W@      @             �H@      [@              @     @S@      @     Pq@      5@      j@      K@       @              7@     �C@      �?      (@      B@      (@     �L@      0@     �T@     �C@       @              @       @               @       @               @       @      @      �?                              �?               @                       @              @      �?                      @      �?                       @                       @                        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?DP�+>i@�	           ��@       	                    �?�4����@�           ��@                          �<@FO��`@9           �@                           �?��A�@           �{@������������������������       ����[o@}             i@������������������������       �d���E@�            �n@                            �?A����@%             O@������������������������       �n#����?             @@������������������������       �{��L^�@             >@
                            �?K�GB�@�           �@                           @���1�Z@g            �e@������������������������       ��sO�=b@A            @]@������������������������       �-o����?&             M@                           �?����<c@Z           ��@������������������������       �罏��# @�            �r@������������������������       ��ߣu�@�             m@                          �7@��j��G@�           �@                           �?�G��X@�           d�@                          �2@t��e�@S             `@������������������������       ��zY .@            �I@������������������������       �Zr(���@4            �S@                          �1@\9��@<           `�@������������������������       �T��k�(@�            �t@������������������������       �S�	���@_           0�@                           @�B5Vv	@$           ��@                          �:@�����$
@h           Ё@������������������������       ���"�	@�             o@������������������������       ����K[
@�            t@                           @Ȫ4�{�@�            �s@������������������������       ��Rf1l�@Q             a@������������������������       �O�[Z	@k             f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        =@     `r@     H�@      ?@     �F@     @~@     @U@     ��@     `k@     ��@     �v@      B@             @R@      e@      @       @      [@      (@     �{@      F@     p@     �V@      @              E@     @V@      @       @      O@      @     @Z@      @@     @X@     �L@       @              D@      T@      @      @     �K@      @     �X@      >@      V@      A@       @              ,@      >@      @      @      9@      @     �G@      5@      <@      4@                      :@      I@              �?      >@              J@      "@      N@      ,@       @               @      "@              @      @              @       @      "@      7@                      �?      @              �?                              �?      @      4@                      �?      @              @      @              @      �?      @      @                      ?@      T@                      G@      @      u@      (@      d@      A@      �?              �?      7@                      "@      @     @U@      @      B@      *@      �?              �?      7@                      @      �?     �G@              ;@      *@      �?                                              @      @      C@      @      "@                              >@     �L@                     �B@      @     `o@      "@      _@      5@                      2@      ?@                      4@              d@      @     �L@       @                      (@      :@                      1@      @     �V@      @     �P@      *@              =@     �k@      v@      8@     �B@     �w@     @R@     �@     �e@     ��@     �p@     �@@      1@     �`@     �n@      *@      8@     �l@     �A@     @}@      V@     �w@     @d@      2@      @       @      9@              @      6@      @      1@      ,@      0@      .@                               @                      @              ,@      @      @      "@              @       @      1@              @      .@      @      @       @      "@      @              *@     �_@     �k@      *@      4@      j@      ?@     0|@     �R@     �v@     `b@      2@      @      1@     �K@              �?      5@      �?     �\@      $@     �R@     �A@              $@     �[@     �d@      *@      3@     �g@      >@      u@      P@      r@      \@      2@      (@     �U@     �Z@      &@      *@      b@      C@     �[@     �U@     �b@     @[@      .@      &@     �L@     �R@      $@      $@     �W@     �A@      J@     �Q@     �O@     �S@      *@              5@      B@       @      @      J@      1@      ;@     �A@      ;@      5@       @      &@      B@     �C@       @      @      E@      2@      9@      B@      B@      M@      @      �?      =@      ?@      �?      @     �I@      @     �M@      0@     �U@      >@       @      �?      &@      @              �?      ;@              :@       @     �A@      4@       @              2@      9@      �?       @      8@      @     �@@       @      J@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��H8hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @>
��@�	           ��@       	                    �?�?ڰ9	@w           V�@                          �<@v�OJ�{@�           0�@                           �?�3m�*@|           X�@������������������������       �e݀�@k            �e@������������������������       ���c��@           �{@                          @@@j�ߡ�@#            �M@������������������������       ��;E�@             F@������������������������       �H�k�qc@	             .@
                          �3@-����	@�           �@                            �?r˟&�B@            z@������������������������       �Y�huU@M             _@������������������������       ������@�            `r@                           @oe�9$
@�           ��@������������������������       ��ο�
@e           �@������������������������       �'�2��{	@c            �d@                           �?7ޛ�%@%           x�@                          �5@'�6�� @a            �@                          �3@�C����?�            Px@������������������������       �����8�?�            �r@������������������������       �O�t�p�?=             W@                            @X���@g            �c@������������������������       �����@S            �`@������������������������       ���b�^�?             ;@                            �?�c8�M@�           �@                           @;�;UL@�           Є@������������������������       �#I���@�            �@������������������������       ��
�)�@             6@                           �?��.,@3            ~@������������������������       �6F;p�@�            �l@������������������������       �p�?P�@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     �q@     �@      G@     �R@     �}@     �T@     ��@     `j@     �@     pu@      B@      7@     �h@      s@     �@@     �N@     �t@     �P@     �w@      e@     0x@     @m@      ?@      �?     �Q@     @S@       @      &@     �V@       @      e@      ?@     `d@      J@      @      �?     �P@     @P@       @      @      T@       @     �d@      9@     `c@     �D@      @      �?      0@      1@                      1@             �I@      @     �M@       @                     �I@      H@       @      @     �O@       @     �\@      6@      X@     �@@      @              @      (@              @      &@              @      @       @      &@                       @      $@                      @              @      @      @      &@                      �?       @              @      @                              @                      6@      `@     `l@      ?@      I@     `n@      M@     @j@      a@      l@     �f@      <@       @      ?@      I@      �?      &@      J@      @      Y@     �F@     �P@      F@      @              @      *@                      4@             �@@      .@      ;@       @      �?       @      8@     �B@      �?      &@      @@      @     �P@      >@      D@      B@      @      ,@     �X@      f@      >@     �C@     �g@     �J@     �[@      W@     �c@     @a@      8@      &@      U@     �b@      <@     �A@      d@      G@     @X@      O@     �b@     �]@      1@      @      ,@      =@       @      @      >@      @      *@      >@       @      3@      @      @     @T@     `j@      *@      ,@     �a@      1@     �@     �E@      z@     @[@      @               @     �S@      @      �?      7@      @     �p@       @     �`@      4@       @              @     �L@              �?      ,@             �j@       @     �V@      @       @              @      ?@                      "@              e@       @     @R@      @       @                      :@              �?      @             �E@              1@                               @      5@      @              "@      @      K@      @      F@      .@                      �?      4@      @               @      @     �A@      @     �C@      .@                      �?      �?                      �?              3@              @                      @     @R@     �`@      "@      *@     �]@      *@     pw@     �A@     �q@     @V@      @             �G@     @S@      @      @     �N@      $@     �j@      7@     �d@     �L@                      E@     @S@      @      @     �N@      @     �j@      4@      d@     �L@                      @              @       @              @       @      @      @                      @      :@      L@      @      @     �L@      @      d@      (@     �]@      @@      @      @      *@      ?@      @      @      =@             @Q@      @     �J@      2@       @              *@      9@              @      <@      @      W@      @     @P@      ,@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ|��0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�(r�l�@�	           ��@       	                   �5@vxs�0@           ��@                           �?��jq�)@�           H�@                           @��U���@           �y@������������������������       ����?��@j            @c@������������������������       �-�I���?�             p@                          �2@��~5A@�            �v@������������������������       ����Y @�            �j@������������������������       ��Y�k%i@`            @c@
                          �9@P���r@-           P~@                            @�7o��D@�            `q@������������������������       �;�A��@m            �f@������������������������       �?iwZa@9            �W@                          �>@ιI$�@�            �i@������������������������       ���_�@i            �d@������������������������       �Kuf��@            �D@                           @lg;�x�@x           ��@                           @|#:z�@�           ��@                          �2@SX��ܮ@�           ��@������������������������       ��&��ۧ@�            pr@������������������������       ��`��7�@�           D�@                          �9@ɰ��|@            �D@������������������������       ���v��@             9@������������������������       �i	\��p@             0@                          �4@ev�L?@�           �@                          �0@?�g@p           ��@������������������������       ��(�[��?&             L@������������������������       ��X�y!�@J            �@                           @3E��$8@e           ��@������������������������       ���SS� @�            x@������������������������       ��S���@r            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �o@     ��@      2@      G@     �}@     �S@     x�@     @i@     X�@     �w@      B@             �R@      g@      @      $@     �X@      @     }@     �E@     0r@     �S@       @              >@     �Y@      �?      @     �J@             �u@      3@      g@      @@      @              4@      G@      �?      @      >@             �g@      0@     �T@      3@                      &@      3@      �?      @      2@              G@      (@     �A@       @                      "@      ;@               @      (@              b@      @     �G@      &@                      $@     �L@              �?      7@             @c@      @     �Y@      *@      @              @      4@              �?      1@             @Y@             �M@       @      @              @     �B@                      @             �J@      @      F@      @                      F@     �T@      @      @      G@      @     @^@      8@     �Z@     �G@      @             �@@     �G@      @              8@             @T@      @     �L@      8@      @              :@      ;@      �?              ,@             �L@      �?     �A@      1@      @              @      4@       @              $@              8@      @      6@      @                      &@     �A@              @      6@      @      D@      4@     �H@      7@                      @      A@              �?      ,@      @      A@      &@     �E@      3@                      @      �?               @       @      �?      @      "@      @      @              *@     @f@     py@      ,@      B@     �w@     �R@     ��@     �c@     @�@     �r@      <@      (@      ^@     �o@       @      :@     �p@     �O@     `h@     �_@      k@     `h@      8@      @     @]@     @o@       @      :@     p@     �O@     `h@      ]@     �j@      h@      3@      �?      5@     �H@              @      E@              P@      8@      K@     �A@       @      @      X@      i@       @      7@     �j@     �O@     ``@      W@      d@     �c@      1@      @      @      @                      "@                      $@       @       @      @       @      @       @                      @                      @               @      @      @              �?                      @                      @       @               @      �?      M@     @c@      @      $@     @\@      &@     �u@     �@@     �r@     �Z@      @              8@     �R@       @      @     �D@       @     �j@      0@     @c@      D@                              @                      �?              >@              0@      @                      8@     �Q@       @      @      D@       @     �f@      0@     @a@     �A@              �?      A@      T@      @      @      R@      "@     �`@      1@     �b@     �P@      @      �?      8@      J@       @             �I@      @      [@      @     @Y@     �@@       @              $@      <@       @      @      5@      @      :@      $@      H@     �@@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ� �NhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@J� YX@�	           ��@       	                    �?j*�?@\           �@                           @0x�)	�@v           X�@                           �?6�~���@�             q@������������������������       �}�z>;@@            �X@������������������������       ���#W;@q            �e@                            @7) ��p@�            �s@������������������������       ��5�4M@o            �d@������������������������       ������@V            �b@
                           @u#2<�
@�           �@                           @*9���@�            0r@������������������������       �x�9@B            �[@������������������������       �Ɔ6uAI@i            �f@                            �? �'U@;           ��@������������������������       �m��m�@M           ��@������������������������       ���J1��@�            @x@                          �<@m���@7           ��@                           �?�O.�B@w           P�@                           �?�$G��	@�           ��@������������������������       ���B\�@�            �i@������������������������       �'ʢ�E
@t           P�@                           �?�(�07@|           ��@������������������������       �_�{��?@�             p@������������������������       ��!�h��@�           ��@                           @�s���	@�            s@                           @D��j	@�            `l@������������������������       ��<�@�            �i@������������������������       ��4F@             4@                            �?4��x@4            �S@������������������������       ���c��4@             C@������������������������       �s�Яq�@             D@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     x�@      =@      N@     �{@     @Y@     ��@      j@     P�@     �x@      7@             �V@      o@       @      2@     �e@      5@     P�@     �R@      x@      c@      @              B@     @R@      @       @     �Y@      *@      `@     �F@     �W@      S@      @              ,@      E@                      @@      @     �R@      4@     �I@     �A@      �?               @      $@                      1@      @      A@      "@      .@       @      �?              (@      @@                      .@              D@      &@      B@      ;@                      6@      ?@      @       @     �Q@      $@      K@      9@      F@     �D@      @              *@      6@      @      @     �@@      @     �@@      2@      .@      4@      �?              "@      "@              @      C@      @      5@      @      =@      5@      @              K@      f@      @      $@     �Q@       @     �~@      =@     0r@     @S@                      &@      K@       @      @      A@      @     @W@      "@      Q@      *@                      @      "@              @      *@             �G@      @      @@                              @     �F@       @      �?      5@      @      G@      @      B@      *@                     �E@     �^@       @      @      B@      @     �x@      4@     �k@      P@                      .@      P@      �?       @      :@             `l@      @     �a@     �F@                      <@      M@      �?      @      $@      @     @e@      *@      T@      3@              0@     �h@     `s@      5@      E@     �p@      T@     �x@     �`@     �x@     �n@      1@      (@     `d@      q@      3@      <@     @m@     �P@     pv@     �Y@     w@     `e@      .@      &@     @X@      a@      1@      4@     �\@      >@     �S@      P@      `@     @T@      &@      �?      :@      A@      �?              @@      �?      7@      @     �M@      2@       @      $@     �Q@     �Y@      0@      4@     �T@      =@     �K@     �L@     �Q@     �O@      "@      �?     �P@      a@       @       @     �]@      B@     �q@      C@      n@     �V@      @              0@      D@                      2@       @      Y@       @      M@      0@              �?      I@     @X@       @       @     @Y@      <@     �f@      B@     �f@     �R@      @      @     �@@      B@       @      ,@     �@@      ,@      B@     �@@      7@     �R@       @      @      9@      8@       @      ,@      5@      *@      .@      ?@      ,@      O@       @      �?      7@      4@       @      ,@      5@      (@      ,@      ;@      ,@      M@      �?      @       @      @                              �?      �?      @              @      �?               @      (@                      (@      �?      5@       @      "@      *@                      @      (@                      @      �?      @              @      @                      @                              "@              ,@       @      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �2@�$6U�@�	           ��@       	                    @0C��@�           <�@                           �?)Q��;i@7           �~@                          �1@|v�7A�@m            `f@������������������������       ��&�R�@A             [@������������������������       ���s�@,            �Q@                            @\���t�@�            `s@������������������������       �`G\�@x             f@������������������������       �C
�{c�@R            �`@
                           @�FwBY� @g           0�@                           �?x7���?           �x@������������������������       �3�����?m            �e@������������������������       �"`��4� @�             l@                           @c'��@c             c@������������������������       ����zC�@E            �Y@������������������������       �i.?� @            �H@                          �;@x/��c@           t�@                           @�ٻ���@�           �@                           �?��bѵ&	@�           x�@������������������������       ��ojO�@�            �x@������������������������       ��(��9�	@�           X�@                           @��^�@m           `�@������������������������       �� ���@c           ��@������������������������       ��t��ѵ@
             5@                           �?�����	@            {@                            @�F����	@�            �p@������������������������       ��6+&�t	@d            �c@������������������������       �� X���	@E            �[@                          @@@ֺ75g@j            �d@������������������������       �(��5�2@[            �a@������������������������       �v��4^@             7@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     r@     0�@      B@     @P@      |@     �V@     ��@     �l@     ��@     `w@     �B@       @      G@     @`@              (@      W@      @      z@     �G@     �k@     �P@      @       @      ;@     �P@              "@     �M@      @     �a@     �E@      X@      C@       @       @      @      4@                      ;@       @     @P@      3@      <@      (@              �?      @      ,@                      (@             �C@      .@      0@      @              �?              @                      .@       @      :@      @      (@      @                      7@      G@              "@      @@      @     @S@      8@      Q@      :@       @               @      9@                      ,@       @     �L@      .@      E@      (@       @              .@      5@              "@      2@      �?      4@      "@      :@      ,@                      3@      P@              @     �@@              q@      @      _@      <@      �?               @     �F@                      1@             �j@      @      X@      ,@                       @      &@                      @             �]@      �?      @@      @                      @      A@                      *@             �W@      @      P@      $@                      &@      3@              @      0@              N@              <@      ,@      �?              $@      .@                      $@              H@              0@      @      �?              �?      @              @      @              (@              (@      &@              &@     `n@     @z@      B@     �J@     @v@     @U@     ��@      g@     ��@     @s@      A@      @     �h@     �u@      =@      E@     �r@     �M@     `�@     `c@     @�@     @m@      ?@      @     @c@     @h@      6@      A@     `j@      E@     �j@      `@      p@     �b@      :@             �M@      G@      @      $@     �D@      �?     @W@      2@     �V@      =@      �?      @     �W@     �b@      2@      8@     @e@     �D@     �^@     �[@      e@     @^@      9@      �?      F@     �b@      @       @     @V@      1@     Ps@      ;@     `p@      U@      @      �?      E@     �b@      @       @     �U@      &@     Ps@      ;@     Pp@     �S@      @               @       @       @              @      @                      �?      @              @     �F@     �R@      @      &@      L@      :@      H@      =@      J@     �R@      @      @      ?@      H@      @       @      =@      3@      5@      5@      5@      K@      @      @      .@      7@      @      @      2@      &@      "@      2@      (@     �C@       @       @      0@      9@      @      @      &@       @      (@      @      "@      .@      �?              ,@      ;@              @      ;@      @      ;@       @      ?@      4@                      *@      6@              @      9@      @      ;@      @      9@      .@                      �?      @                       @      @              �?      @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�Y�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?^kj�il@�	           ��@       	                   �;@p1ɇ>W	@           h�@                          �2@Vz�y	@i           p�@                           @Ӳ���@�            �s@������������������������       ����P�@�            �n@������������������������       ����}[@,             Q@                          �:@d:ҫ�y	@�           ��@������������������������       ��P��s	@v           ؎@������������������������       ��#�.a�@)            @R@
                          �<@��-k	@�            �o@                           �?4�@�@$             L@������������������������       ��U��@
             .@������������������������       �Q��-gx@            �D@                           @h4Sb�;	@�            �h@������������������������       �T�
�=F@x             f@������������������������       ��tR~�E@             5@                          �4@�\q�@�           ޡ@                           @����@�           �@                          �1@v��晩@;            @������������������������       ��B�q=@l            @e@������������������������       �8�5���@�            `t@                           @�iZ+!o@�           ��@������������������������       ��E�l��?#            |@������������������������       ��&��@�             q@                           �?c��|��@�           ��@                          �=@0U@�            �p@������������������������       �r@��\@�            `o@������������������������       ��:�le@
             ,@                          �<@�&�qp@�           �@������������������������       ��SCw1@�           ��@������������������������       ��(p��@<            �X@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@     u@     �~@      9@      J@     0|@     �S@     �@     �k@     `�@     �x@      @@      8@     `h@     �j@      3@      >@      l@     �G@     @j@      b@     �q@     �i@      8@      .@     @d@     �e@      *@      :@     @i@     �B@     @h@     �^@      p@     �b@      5@       @     �C@     �B@               @     �L@      @     �O@      .@     �L@     �A@       @              9@      <@               @     �E@             �M@      "@     �I@      ;@               @      ,@      "@                      ,@      @      @      @      @       @       @      *@     �^@     @a@      *@      8@      b@      A@     ``@     �Z@     �h@     �\@      3@       @     @^@     �`@      *@      8@     @`@     �@@     @]@     @Y@     `g@     �Y@      3@      @       @      @                      .@      �?      ,@      @      (@      (@              "@     �@@      D@      @      @      7@      $@      0@      7@      =@      M@      @      @      &@      $@               @      @      @      @              @      &@               @              �?                      @              �?              @      @               @      &@      "@               @      �?      @      @              @      @              @      6@      >@      @       @      2@      @      (@      7@      7@     �G@      @       @      4@      ;@      @       @      0@      @      &@      1@      6@     �G@              @       @      @                       @              �?      @      �?              @       @     �a@     0q@      @      6@     @l@      ?@     x�@     �S@     x�@     `g@       @              P@     `a@      �?      *@     �T@      @     �@      B@     0r@      R@      �?             �B@     �Q@              @     �G@      @     @g@      8@     �U@     �B@                      @      5@                       @             @U@       @      ?@      (@                      @@     �H@              @     �C@      @     @Y@      0@     �K@      9@                      ;@     @Q@      �?       @      B@       @     �t@      (@     �i@     �A@      �?              $@      C@              �?      (@             @l@      @     �a@      2@                      1@      ?@      �?      @      8@       @     �Y@      @     @P@      1@      �?       @     �S@      a@      @      "@     �a@      9@     �p@      E@     �m@     �\@      @              *@      A@                      5@      @     �[@      @      N@      0@       @              *@     �@@                      4@      @      [@      @      M@      &@                              �?                      �?               @      �?       @      @       @       @     @P@     �Y@      @      "@     �^@      6@     �c@      B@      f@     �X@      @       @      J@     �V@      @      @     �W@      3@     �b@      @@      e@     �S@      @              *@      &@              @      <@      @      "@      @       @      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJA��;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?t�@�	           ��@       	                    �?&��"2@'           �@                            �?��:�|�@2           `~@                          �5@~�1e��@W             a@������������������������       ����@'            �O@������������������������       �W!h`A@0            �R@                          �<@�|����@�            �u@������������������������       ����dT@�            �r@������������������������       �=��Y��@            �J@
                          �>@���g�@�           ��@                           �?q� /v@�           @�@������������������������       �����@           �|@������������������������       �<�rl�@�            �s@������������������������       ���Dh�@             4@                          �1@��l	D"@�           ��@                          �0@����vY@�            �u@                           @��V�@G            @W@������������������������       �b��Ѐ�@!            �F@������������������������       �Wd�ګ�?&             H@                           @	�4+.@�             p@������������������������       �`0d���?             B@������������������������       ��8�B@�            �k@                           @��;b̏@�           С@                          �;@4{_S	@�           D�@������������������������       �雍L��@S           D�@������������������������       ��0�c	@�             p@                           @�e��d@�           ��@������������������������       �H�:6@            {@������������������������       ���M@�            pr@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        =@     �q@     ��@      7@      H@     �}@     �Q@     �@     @i@     @�@     pv@      >@              T@     �g@      @      @     �\@       @     p|@      C@      s@     @T@      @             �H@      T@      @      @      M@      @      X@      8@     �]@      G@      �?              0@      =@                      2@       @      8@      @      ?@      *@                              0@                      @              0@      �?      2@      @                      0@      *@                      (@       @       @      @      *@      @                     �@@     �I@      @      @      D@       @      R@      4@      V@     �@@      �?              >@     �F@      @       @      >@       @     �Q@      1@     �S@      0@      �?              @      @              @      $@              �?      @      $@      1@                      ?@      [@               @      L@      @     pv@      ,@      g@     �A@       @              >@     @Z@               @     �J@       @     0v@      $@      g@      @@       @              3@      Q@               @      B@      �?     �l@      @     �T@      2@                      &@     �B@                      1@      �?     �_@      @     �Y@      ,@       @              �?      @                      @       @      @      @              @              =@     �i@     `w@      3@     �D@     `v@      O@     ؁@     �d@     �@     `q@      ;@              .@      E@      �?       @      6@      �?     �a@      1@     �T@      ;@                      @      .@                      @             �@@      �?      5@      (@                      @      (@                      @               @      �?      @      @                              @                                      9@              .@      @                      &@      ;@      �?       @      .@      �?      [@      0@      O@      .@                       @                                              6@      @       @      @                      "@      ;@      �?       @      .@      �?     �U@      $@      N@      &@              =@     �g@     �t@      2@     �C@      u@     �N@     �z@     `b@     Pz@     `o@      ;@      =@     `b@     �m@      (@      =@     �o@     �I@     @m@     �`@     �j@     �g@      8@      2@     �_@     �j@      "@      ;@      k@      B@     �k@     @[@     �e@     ``@      1@      &@      5@      7@      @       @      B@      .@      ,@      8@     �D@     �M@      @              E@     �W@      @      $@     �T@      $@     �h@      ,@     �i@     �N@      @              2@      L@      �?      �?      G@             �a@      &@     �_@      =@                      8@     �C@      @      "@     �B@      $@     �J@      @      T@      @@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�=AhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ni]�@~	           ��@       	                   �5@���DV�@�           T�@                          �1@��y�@�           P�@                           �?`�&dP��?�            �n@������������������������       ��Qc�6�?O            �_@������������������������       ��9LnU��?L             ^@                           @�\��<�@*           0}@������������������������       �]H�$^r@�            `m@������������������������       �.[���?�             m@
                          �<@8�>�q�@           �|@                            @� ' �@�             w@������������������������       �h�n@�            0p@������������������������       �+3��j@F            �[@                            @>�{3��@8            @V@������������������������       ��Pn-�@*             P@������������������������       �0R\�@             9@                          �5@�0��@�           h�@                           @��\�u�@�           ��@                           @ס��ߔ@K            �@������������������������       �,�x��@4           �}@������������������������       ��uǰ]@            ~@                           @�m�z@H           X�@������������������������       �آ���@4           @�@������������������������       � W�n 	@            �A@                          �;@��l
�@           $�@                           @��]��@=           X�@������������������������       ����N@�           @�@������������������������       ��W\XV@T            ``@                          @@@��P	��@�            �s@������������������������       �Y%�
�)	@�            q@������������������������       ��5��:�@            �F@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     @�@      6@      Q@     �y@     �R@     Ȑ@     @j@     ��@     @t@      ?@             @U@     �b@       @      ,@     @S@      (@      }@      A@     �p@      Q@      @             �F@     �U@      �?      @      >@      @     �u@      0@     �b@      =@                      @      ;@               @      $@              b@      @      G@      $@                       @      .@               @      @             �R@       @      0@      "@                       @      (@                      @             �Q@      �?      >@      �?                     �D@     �M@      �?      @      4@      @     �i@      *@     �Y@      3@                     �@@      =@      �?       @      0@      @     @R@      &@      J@      ,@                       @      >@              �?      @             �`@       @      I@      @                      D@     �O@      �?      "@     �G@       @     �\@      2@      ]@     �C@      @             �A@     �I@      �?      @      @@       @     �X@      (@      Z@      8@       @              <@      @@      �?              9@       @     �O@      @      S@      4@       @              @      3@              @      @             �A@       @      <@      @                      @      (@              @      .@              0@      @      (@      .@       @              @      &@               @      @              (@      @      (@      ,@       @              �?      �?              @      (@              @       @              �?              ,@     �l@     0y@      4@      K@      u@     �O@     �@      f@     H�@      p@      ;@      $@     �T@      l@      $@      9@      e@      0@     �z@     @R@     �u@     @\@      0@      @     �I@     �a@       @      &@      [@      "@     �p@      ?@     �o@     �S@      �?      @      A@     �P@      @      "@     @Q@      @     @W@      :@     �Z@     �K@      �?              1@     �R@      �?       @     �C@       @     �e@      @     @b@      7@              @      @@      U@       @      ,@      N@      @     �d@      E@      W@     �A@      .@              ?@      S@       @      &@      L@      @     �d@     �D@     �U@     �@@      *@      @      �?       @              @      @      �?       @      �?      @       @       @      @      b@     @f@      $@      =@      e@     �G@     `f@     �Y@      j@     �a@      &@      �?     �Z@     �a@      @      8@     �]@      =@     �b@     @T@     `d@     �S@      "@             @T@     �]@      @      8@     �Z@      9@     ``@      M@      c@      R@      @      �?      9@      6@       @              (@      @      4@      7@      &@      @      @      @     �C@      C@      @      @      I@      2@      <@      6@     �F@     @P@       @      @     �@@      ;@      @      @      G@      2@      ;@      4@      C@     �I@       @              @      &@                      @              �?       @      @      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?t��>�@�	           ��@       	                    �?��^��n	@           P�@                           �?���I�@�           ��@                           �?��	+�@�             o@������������������������       ��}���a@9            @V@������������������������       ���s�@f            �c@                           �?~�ef�@�            pv@������������������������       �q���@B             Z@������������������������       ���#��@�            �o@
                          �;@�ɘ�_�	@�           ��@                           �?YI�Z�	@           ��@������������������������       �bc��T�	@�            �r@������������������������       �f��I	@J           X�@                           @4l��	@z            @h@������������������������       ������@T            �_@������������������������       �Vm��^�@&            �P@                           �?��q @�           �@                          �2@�Ĭ�@�           ��@                            @f��  @�            �r@������������������������       �@�$� @�            �m@������������������������       ����H�?&            �M@                            @����@            {@������������������������       ����6n@�            @v@������������������������       ���=�@2            �S@                           @�����@@�           d�@                           @����Ii@           �{@������������������������       �S�󔖝@�            �q@������������������������       ����d@a            �c@                           @(Bk�A@�           t�@������������������������       ��,�o��@�            �@������������������������       ��zCH�~@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     pr@     ��@     �B@     �N@     �{@     @U@     �@     �n@     �@     �w@      4@      6@     �g@     �m@      7@      C@     �k@      J@      k@      d@     �o@      h@      ,@       @     �B@     @[@      @      "@      T@      $@     �^@      G@     @]@     �P@      @      �?      7@      G@      �?      �?      F@      @      L@      .@     �B@      3@      �?               @      &@                      "@             �@@      �?      8@      @              �?      .@     �A@      �?      �?     �A@      @      7@      ,@      *@      0@      �?      �?      ,@     �O@       @       @      B@      @     �P@      ?@      T@     �G@      @              "@      6@                      @              :@       @      @@      @       @      �?      @     �D@       @       @      >@      @     �D@      =@      H@      E@       @      4@     �b@     �_@      4@      =@     �a@      E@     �W@     �\@     @a@     �_@      "@      (@      _@     @Z@      ,@      5@      `@      :@      U@      W@     �]@     �U@      "@       @     �F@      B@      "@      @     �A@      ,@      >@      F@      @@      E@      �?      $@     �S@     @Q@      @      .@     @W@      (@      K@      H@     �U@      F@       @       @      ;@      6@      @       @      ,@      0@      $@      6@      4@     �D@              @      0@      6@      @      @      @       @       @      "@      0@      ?@              �?      &@                      @       @       @       @      *@      @      $@                     �Z@     `t@      ,@      7@      l@     �@@     P�@     @U@     �@     @g@      @             �@@     �V@      �?      �?     �H@      @     @u@      &@     �d@      C@                      $@     �A@                      4@             �c@              K@      6@                      "@      ?@                      3@             �]@             �D@      4@                      �?      @                      �?              C@              *@       @                      7@     �K@      �?      �?      =@      @     �f@      &@     �[@      0@                      3@      I@      �?              5@      @      c@      &@     �U@      &@                      @      @              �?       @              ?@              8@      @                     �R@     �m@      *@      6@      f@      <@     `{@     �R@     �u@     �b@      @              7@     @U@              $@      N@      *@     �W@      H@      N@      I@      �?              .@     �J@              @     �E@      &@     �I@      6@     �D@     �E@      �?               @      @@              @      1@       @     �E@      :@      3@      @                     �I@     �b@      *@      (@      ]@      .@     �u@      :@     �q@     �X@      @              ?@     �[@      @       @     �R@      @     q@      1@     �h@      L@      @              4@      D@      $@      $@      E@      (@     �Q@      "@      V@      E@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$�:hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �;@��/AX@�	           ��@       	                   �1@0��y��@�           ��@                           �?g���@�           ��@                           �? @��ϕ@�            Ps@������������������������       ��s��_��?S             a@������������������������       ��/��@i            �e@                            @}���]@�            �s@������������������������       �ġH�@�            �l@������������������������       ��o�m@8             V@
                          �8@C(�R@           �@                           @��6�@�           h�@������������������������       ���Z<j�@*           �@������������������������       �-�&X��@�           ��@                           @��'@�A@4           @}@������������������������       �v��;@           �y@������������������������       �&8(m�-@"            �K@                           @ȇ�W��	@            �|@                           @�h`$��	@�            �p@                           �?6>p7�	@            �h@������������������������       ��l�p�@:            @X@������������������������       ���Bq
@E            @Y@                           �?T���M@)            �P@������������������������       �V�Џ�@            �C@������������������������       ��;���@             ;@                           @ -�ե�@x            �h@                           �?�P���@(            �P@������������������������       �t�͊�:@             ;@������������������������       �TL�x8@             D@                          @@@<<�ɞG@P            @`@������������������������       �+r|6F�@E            @\@������������������������       �)���	@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �s@     ��@     �@@      N@     `y@      U@     ��@      m@     h�@     �u@      ;@      @     �p@     �@      9@     �H@     u@      O@     P�@      h@     x�@     pp@      7@      �?      B@      R@      �?      @     �A@             �q@      6@     @a@      C@              �?      ,@      @@      �?      @      4@             @b@       @      L@      <@                      @      .@                      *@             �S@       @      0@       @              �?      $@      1@      �?      @      @              Q@      @      D@      4@                      6@      D@              �?      .@             �`@      ,@     �T@      $@                      *@      ;@                      *@             �X@      (@     �O@      @                      "@      *@              �?       @             �B@       @      3@      @              @     �l@      {@      8@     �F@     �r@      O@     ��@     `e@     (�@      l@      7@      @     �g@     �w@      2@      B@      o@      I@     ��@     �[@      �@     �g@      3@      @     ``@     �i@      (@      ?@     �e@      B@     �k@     @X@     �n@     �\@      .@             �M@     �e@      @      @     @S@      ,@     `w@      *@      q@     �R@      @      �?      D@     �K@      @      "@     �J@      (@     @W@     �N@     @X@     �B@      @              <@      I@      @      "@     �I@      (@     �S@      I@     �V@      B@      @      �?      (@      @       @               @              ,@      &@      @      �?      �?      $@     �J@     �L@       @      &@     @Q@      6@     �C@      D@      O@     �U@      @      "@      8@      C@       @      @      >@      ,@      ?@      1@      C@      J@      @      "@      6@      <@       @      @      ;@      (@      *@      $@      <@      D@      @      �?      3@      &@               @      (@       @      @      @      2@      5@               @      @      1@       @       @      .@      $@      @      @      $@      3@      @               @      $@               @      @       @      2@      @      $@      (@                       @      "@              �?      �?      �?      .@               @       @                              �?              �?       @      �?      @      @       @      $@              �?      =@      3@      @      @     �C@       @       @      7@      8@      A@      �?               @      @      @      @      5@       @              @      @      "@                      @      @       @      �?      $@                      �?              @                      @      �?      @       @      &@       @              @      @      @              �?      5@      (@               @      2@      @       @      0@      4@      9@      �?              3@      @               @      .@      @       @      0@      3@      6@      �?      �?       @      @                      @                              �?      @        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��L(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?P�C�>:@�	           ��@       	                    @`����@
           \�@                          �<@�z����@�           ��@                            �?U%��@@{           P�@������������������������       ���C�k$@�            `u@������������������������       �WJ�@�            @q@                           �?n!��@4            @S@������������������������       �,>K(�, @
             0@������������������������       �豀�Zi@*            �N@
                           �?ó
��� @[            �@                            �?�P��,= @�            �s@������������������������       ����B<�?(            �L@������������������������       ��ؓ� @�            �o@                           @k���a� @�             m@������������������������       ���8�|�?X            �a@������������������������       �^���ۜ@9            @V@                          �4@h�Fo@�           �@                          �1@�Ab?�@�           L�@                           �?����Z�@�            pv@������������������������       �q=�B�}@p            �f@������������������������       �,~�J�x@j            `f@                           @g�	�~�@           `�@������������������������       �Y��G>�@�            �w@������������������������       ��/I��,@           0{@                           @�1r��@�           |�@                           �?r<ͤ��@�           ��@������������������������       ��N�}�K	@F            �\@������������������������       ���D���@I           Ԕ@                           @4��o@"             L@������������������������       ��i��V�@            �F@������������������������       ��)���?             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �t@      �@      7@     �K@     0|@     �T@     ��@     �m@     �@     �t@      ?@      �?     �W@     �f@      @      ,@     @Z@      &@     �z@     �F@     �q@     �P@      @      �?      S@      [@      @      &@     �R@      @     �d@      C@     `c@     �J@      @      �?     @P@     @X@      @      @     �P@      @      d@      <@      b@      A@      @      �?      @@     �K@      @       @      >@       @     �U@      3@      V@      3@      @             �@@      E@      �?      @      B@      @     �R@      "@     �L@      .@                      &@      &@              @       @              @      $@      $@      3@      �?              @      @                                       @              �?       @                      @      @              @       @              �?      $@      "@      1@      �?              2@     @R@              @      ?@      @     �p@      @      `@      ,@                      @     �C@              @      ;@      �?      d@      �?      P@      "@                              @                      @              B@              "@      @                      @      B@              @      7@      �?     @_@      �?     �K@      @                      &@      A@                      @      @      Z@      @      P@      @                      @      4@                      �?      @      R@             �C@      �?                      @      ,@                      @              @@      @      9@      @              &@     `m@     �v@      3@     �D@     �u@     �Q@     H�@      h@     8�@     `p@      :@       @      S@     @b@      @      "@     �\@      5@     `w@     �Q@     �n@     @Y@      @      �?      .@      C@      �?       @      ;@      �?      a@      6@      W@      8@              �?       @      3@      �?      �?      1@      �?     @R@      *@      @@      ,@                      @      3@              �?      $@             �O@      "@      N@      $@              �?     �N@      [@      @      @     �U@      4@     �m@      H@     `c@     @S@      @      �?     �A@      J@      �?      @      C@      &@     @]@      (@     �S@      =@                      :@      L@      @      @     �H@      "@     @^@      B@     @S@      H@      @      "@     �c@     �k@      *@      @@      m@      I@     `j@     �^@      q@      d@      5@      @     @b@     `k@      *@      @@     �k@      H@      j@     @Z@     �p@      d@      3@      @      5@      &@              @      0@      @      @      *@      1@      1@      @      @     @_@      j@      *@      =@     �i@     �E@     �i@      W@     @o@      b@      .@      @      *@       @                      $@       @       @      1@      @               @      @      @      �?                      "@      �?              1@      @               @              @      �?                      �?      �?       @                                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJD�oqhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?n��O�@�	           ��@       	                    @F>,���@           ��@                           �?/�/��@�           X�@                          �8@���A@�            pt@������������������������       �Ɗ��@�            �k@������������������������       �a��J+@>            �Z@                           �?C�JT��@�            @t@������������������������       ���\�2@�            �n@������������������������       �O���ɴ@4            @S@
                           �?09���@p           ��@                            @z�Zk%�@�            �u@������������������������       �>��~#@�            r@������������������������       �*��e\��?!            �N@                           @�L��}R@�            @o@������������������������       �]����?P            �`@������������������������       ��z��|A@I            �\@                            @�y�+=n@�           ̤@                           @�X{��@�           �@                           �?
U�u�t	@L           ��@������������������������       ���m���@�            `q@������������������������       �]�n�	@�           ��@                           @!��]A@U           ��@������������������������       ��A����@�           x�@������������������������       ��6�m�4@�            @p@                           �?뚃�(^	@�           ��@                           �?�<~�St@/             S@������������������������       �I%l�}�@             8@������������������������       ���6�.@!             J@                          �9@�R2e(	@�           ��@������������������������       ����F�@W            �@������������������������       ��$�q��
@i            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     @s@     ��@      ?@     �P@     �|@     @Z@     ��@     �i@     (�@     �v@      ?@      �?     @W@     �d@      @       @     �[@      .@     �z@      D@     �q@     �V@      @      �?     @R@      T@       @      @     �S@      @     �c@      ?@     @b@     �N@      @      �?      @@      D@       @      @      D@      @     �V@      3@      K@      B@      �?              7@      :@       @      �?      ;@      @     �S@      $@     �@@      0@      �?      �?      "@      ,@              @      *@      @      (@      "@      5@      4@                     �D@      D@               @      C@             @Q@      (@      W@      9@      @             �B@      B@               @      ?@             �E@      (@      P@      2@      @              @      @                      @              :@              <@      @      �?              4@     �U@      �?      �?      @@       @      q@      "@     �a@      >@                      *@     �H@              �?      8@      @     �c@      @     �S@      1@                      &@     �G@                      7@      @      `@      @      M@      *@                       @       @              �?      �?              >@              5@      @                      @     �B@      �?               @       @     �\@      @      O@      *@                      @      0@                      @       @     �Q@              B@      �?                              5@      �?              @              F@      @      :@      (@              3@     �j@      w@      <@     �M@     �u@     �V@     x�@     �d@     `~@     �p@      9@      "@     �a@     `p@      0@      D@      m@     �K@      |@      ]@      v@     `f@      *@      "@     �T@     �a@      "@      7@     �b@     �F@     @^@     �U@      `@     �[@      &@              2@      H@      �?      @      G@       @     �H@      0@     �B@      G@      @      "@      P@     @W@       @      3@     �Y@     �B@      R@     �Q@      W@      P@      @             �M@     @^@      @      1@     �T@      $@     pt@      =@     �k@     @Q@       @              D@     @W@       @      @      J@      @      q@      1@     �b@     �G@      �?              3@      <@      @      (@      ?@      @     �K@      (@      R@      6@      �?      $@     �R@     �Z@      (@      3@     �\@     �A@     �a@      H@     �`@     �V@      (@               @      ,@              @      "@      @      �?      .@      @      $@       @                      "@                      �?      @               @              @       @               @      @              @       @       @      �?      *@      @      @              $@     �P@      W@      (@      ,@     �Z@      >@     �a@     �@@     �_@     @T@      $@      @     �G@      T@      @       @     @U@      (@     �]@      7@     �Z@     �I@      @      @      3@      (@      @      @      5@      2@      8@      $@      5@      >@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�d�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�G�B`@�	           ��@       	                   �<@� c��i@�           ��@                            �?�/p��@�           4�@                           �?�0�{t*@u           ��@������������������������       ���S1��@�            �t@������������������������       �ٳ�kb@�            pp@                            @,�߭E@B           �@������������������������       ���\�Ӂ@�            �i@������������������������       ��$�ox�@�            �r@
                           @���L@:            �V@                            �?i"��@*             P@������������������������       �+�C@g�@             A@������������������������       ��Wȹ@             >@                           �? ���@             ;@������������������������       �騼����?             ,@������������������������       ����\a� @             *@                           @oAA0I@�           B�@                           @���2.�@�           ��@                            @Ъ٫�7	@I            �@������������������������       �J��s	@�           Ј@������������������������       �E��;	@S           0�@                           �?.��}��@t            �@������������������������       ��I���/@.             U@������������������������       �3�B�G@F           `�@                           @`+L}�	@�            v@                            �?�{�[P	@|            �i@������������������������       �=�<�@M            @_@������������������������       �����W@/             T@                            �?��ַ��@\            �b@������������������������       ��)\�C@             B@������������������������       �l��6�4@G             \@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        <@     �q@     x�@      9@      N@     �|@     �U@     ��@     �l@     ��@     pu@      >@             �R@     �c@       @      *@     �Y@      *@     �{@      F@     q@     �P@      @             @Q@     �a@       @      $@     @V@      &@     �z@     �A@     �p@     �H@      @              E@     �T@       @      @      J@      @     �j@      *@     �b@      9@      @              :@      D@      �?      @      ?@      @     @`@      (@      O@      0@       @              0@     �E@      �?              5@             �T@      �?      V@      "@       @              ;@     �M@              @     �B@      @     �j@      6@     �\@      8@                      &@      6@                      &@      @     @W@      (@      F@      @                      0@     �B@              @      :@       @      ^@      $@     �Q@      1@                      @      1@              @      ,@       @      0@      "@       @      1@                      @      *@              @      &@              @      "@       @      0@                      @      @               @      @               @      @       @      ,@                       @      $@              �?      @              @      @               @                              @                      @       @      &@              @      �?                              @                               @       @              �?                                      �?                      @              @              @      �?              <@     �i@      y@      7@     �G@     Pv@     �R@     ��@      g@     h�@     Pq@      :@      2@     �e@     �u@      5@     �F@     �s@     �K@     (�@     �a@     0~@      n@      .@      0@     �^@     �h@      3@      >@     �k@     �C@      h@     @]@     `j@     @d@      .@      "@     �R@      V@      @      8@     �`@      8@     �]@     �S@     �`@     @X@      @      @      H@     �[@      ,@      @     @V@      .@     �R@      C@      S@     @P@       @       @     �J@     @b@       @      .@     �V@      0@     @t@      8@      q@     �S@               @      @      1@              �?      @      @      .@      @      5@      @                      I@      `@       @      ,@     @U@      "@     Ps@      1@     `o@     �R@              $@      ?@      L@       @       @      F@      3@     �L@     �E@      E@      B@      &@      $@      &@     �C@              �?      =@      0@      1@     �A@      6@      3@      @      @      $@      4@                      1@      (@      @      :@      0@      (@      @      @      �?      3@              �?      (@      @      ,@      "@      @      @       @              4@      1@       @      �?      .@      @      D@       @      4@      1@      @              @      @      �?      �?                      $@      @       @       @                      0@      (@      �?              .@      @      >@      @      2@      "@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJr�!ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?e`DX�k@�	           ��@       	                   �4@��X%�@           8�@                           @b#� �@�           p�@                           �?00Ԅ�@�            �r@������������������������       �.JB@I            �`@������������������������       ����T�A@m             e@                            �?�����?�             v@������������������������       �9c��u��?8             W@������������������������       ���E�� @�            `p@
                          �<@�w�m@r            �@                          �9@�M����@<           p@������������������������       �HQh@x�@�            px@������������������������       �� 4�9@J             \@                          @@@[Ͷ_@6            @R@������������������������       ��9�q`�@'             K@������������������������       ��qI4��@             3@                            @��M@�           ��@                          �6@ 'e���@�           L�@                           @o^�Z|u@�           H�@������������������������       ��q̿�3@\           ��@������������������������       ��|2ji@�           ��@                           �?��<`3!	@�           �@������������������������       �m���k@             G@������������������������       ��3}r1�@�           ��@                           �?X��MC	@           @�@                           �?�D��
@4           �}@������������������������       �����m@a             b@������������������������       �I	a�[
@�            �t@                           @~K3��@@�            �t@������������������������       ����}@�            �r@������������������������       �Õ��P�@             B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     0t@     �@      ?@      L@     �|@     @T@     Џ@      j@     (�@     �v@      ?@             @Y@     �d@      @      $@     �Y@       @      {@     �B@      q@     �U@      @              D@     �U@               @     �B@      �?      r@      2@     `a@     �C@      @              8@      B@                      ?@      �?     @X@      (@      R@      9@       @              "@      1@                      5@      �?      G@      @      2@      &@       @              .@      3@                      $@             �I@      @      K@      ,@                      0@     �I@               @      @             �g@      @     �P@      ,@      �?                      0@                                     �I@              5@      @                      0@     �A@               @      @             �a@      @      G@      $@      �?             �N@      T@      @       @     @P@      @     @b@      3@     �`@     �G@       @              I@     �R@      @      @     �K@      @      a@      *@     �_@      =@                     �E@      J@      @      @      D@      @      [@      &@      X@      :@                      @      6@                      .@      @      <@       @      ?@      @                      &@      @               @      $@              $@      @       @      2@       @               @      @                      @              $@      @      @      0@       @              @       @               @      @                       @      @       @              9@     �k@     �w@      9@      G@     0v@     @R@     @�@     �e@     0@     `q@      :@      @     @c@      o@       @     �B@      n@      J@     �{@     �^@     pv@     �g@      .@       @      U@     �b@      @      7@     @a@      3@      v@      L@      m@     @Y@      @              C@     �N@      @      @      G@      &@     �e@      *@     @`@     �I@               @      G@     �V@              0@      W@       @     �f@     �E@     �Y@      I@      @      @     �Q@     @X@      @      ,@     �Y@     �@@      V@     �P@     �_@      V@       @       @      @      @              @      @      �?      �?       @       @      @              @     �O@     �W@      @      @     �X@      @@     �U@     �M@     �]@      U@       @      2@      Q@     @`@      1@      "@     �\@      5@     �a@     �H@     �a@     @V@      &@      2@     �H@     @P@      &@      @     �T@      3@     �K@      A@     �Q@      L@      "@      �?      &@      2@       @      �?      <@      @      <@      $@      4@      3@       @      1@      C@     �G@      "@      @      K@      ,@      ;@      8@      I@     �B@      @              3@     @P@      @      @      @@       @     �U@      .@     �Q@     �@@       @              ,@      L@      @      @      9@       @     �T@      *@     �P@     �@@                      @      "@      @              @              @       @      @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�,hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�Iq:E}@�	           ��@       	                    @<��Љ7@�           L�@                          �2@�����@d           ��@                           @^?	IG@�            �r@������������������������       ���ތ��@�             j@������������������������       �<����k@6            �U@                           �?)B8cj	@�           @�@������������������������       �s/ � @�            �s@������������������������       �9Y��	@�           ��@
                           @�"4�u@�           ��@                           �?i�yT&�@�           Đ@������������������������       �^�W�`�@:           �@������������������������       ���ap��@d           ��@                           @�b���;@�            �w@������������������������       ���"촔@�            Pv@������������������������       �E�2��@             8@                           @V�@= @�           ��@                           �?~���@�           ��@                          �5@D���@�            �i@������������������������       �e���'�@O            �]@������������������������       �A���Y@7            �U@                           �?+ьZLR	@v            �@������������������������       �sJ6��@$             M@������������������������       ����'	@R           P�@                           @4>���Y@�             q@                           @U�-@�            �i@������������������������       ��{F�k��?Q             `@������������������������       ��V��@7            �S@                           6@6i�zAw@'            �P@������������������������       �<��i�x @             @@������������������������       ���P;@            �A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �t@     ��@      ?@     @P@     �|@     @Q@     ��@     �k@     Ј@     x@      <@      $@     �m@     �z@      1@      G@     �s@      H@     8�@      d@     p�@     `q@      2@      $@     �c@     �h@      &@      <@     �h@     �D@     �k@      ]@     @m@      e@      0@              1@      F@                      C@              U@      6@     �L@      A@                      &@      >@                      ;@              P@      @     �I@      7@                      @      ,@                      &@              4@      3@      @      &@              $@     �a@      c@      &@      <@      d@     �D@      a@     �W@      f@     �`@      0@              I@      A@              @      D@      @      O@      ,@     @Q@     �B@       @      $@      W@     �]@      &@      5@     @^@     �B@     �R@      T@      [@     �X@      ,@              T@     `l@      @      2@     @\@      @     �~@     �F@     @v@     @[@       @              C@     `e@      @      1@     �S@      @      w@      @@      r@     �Q@                      .@     �U@      @      @      =@      @      i@      *@     �`@      8@                      7@     @U@       @      ,@     �H@      @      e@      3@     @c@      G@                      E@      L@      �?      �?     �A@      �?     �^@      *@      Q@     �C@       @              @@      L@                     �@@             �]@      (@     �P@     �B@       @              $@              �?      �?       @      �?      @      �?       @       @               @     @W@      b@      ,@      3@      b@      5@     @m@      N@     �i@     �Z@      $@       @     @S@     �_@      "@      .@     �_@      2@     @^@      J@      `@     �W@      $@              2@      :@              @      8@      �?     �I@      @     �H@      :@                      "@       @                      &@      �?      D@      @      =@      1@                      "@      2@              @      *@              &@      @      4@      "@               @     �M@      Y@      "@      &@     �Y@      1@     �Q@      G@     �S@      Q@      $@      @      @      0@               @      ,@       @              "@       @      @       @      @      K@      U@      "@      "@     @V@      .@     �Q@     �B@     @S@     @P@       @              0@      2@      @      @      2@      @     @\@       @      S@      *@                      $@      .@               @      &@              W@       @     �O@      @                      @      "@                      "@              J@      @      I@                              @      @               @       @              D@      @      *@      @                      @      @      @       @      @      @      5@              *@      @                      �?               @              @      @      .@               @                              @      @      @       @      @              @              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ.VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�xujE@�	           ��@       	                    �?�`��@t           `�@                          �;@���D�(@�           ��@                           �?�7�B�Z@_           ��@������������������������       ��gm,�/@�            `x@������������������������       �!���f�@b             c@                            �?o��u�@4            @T@������������������������       �e(ĝ�@            �E@������������������������       ���#���@             C@
                           @����e	@�            �@                           �?L�G�x2	@r            �@������������������������       �X���'x	@�           ��@������������������������       �Ğf��@�            �r@                          �:@/:8�C	@o            �@������������������������       �p�Wb��@            P|@������������������������       �Y}D:v	@O            �^@                          �7@M��o@4           d�@                          �1@�W����@0           ԓ@                           @O).d��?�            �u@������������������������       ���sj=��?u            `f@������������������������       ���@<� @g            �d@                          �4@�Ģ�@T           ،@������������������������       ��o�}��@`           �@������������������������       �X��N�H@�            �w@                          �=@�xE�o�@           @z@                            @c�x%k @�            �u@������������������������       �l�.@�             r@������������������������       �����@)             N@                            �?"!d8@(             R@������������������������       �'*�ED� @             1@������������������������       ����%(@             �K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     x�@      7@      M@     �|@     @W@     (�@      k@     ��@     @v@      =@      1@     �i@     t@      3@      E@     �s@     @R@     x@     @f@     px@     `o@      8@      �?     �K@     �Q@      �?      "@     �S@      @     �d@      ?@      b@     �N@      �?             �G@      O@      �?      @      O@      @     �d@      7@      `@      G@                      A@     �J@      �?      @      J@      @     @W@      6@      W@     �A@                      *@      "@              �?      $@      �?     �Q@      �?      B@      &@              �?       @      "@              @      0@      �?       @       @      1@      .@      �?      �?      @      @                      @      �?      �?      @       @      *@      �?              @      @              @      (@              �?       @      "@       @              0@     �b@     @o@      2@     �@@      n@      Q@     `k@     `b@     �n@     �g@      7@      &@     @X@     ``@      $@      6@     `c@     �H@     �a@      T@     �e@      b@       @      &@     �R@     �V@      $@      2@     @]@      B@     �V@      F@     �_@     �Y@       @              7@      D@              @      C@      *@     �J@      B@     �G@     �E@              @      J@     �]@       @      &@     �U@      3@      S@     �P@     @R@     �F@      .@       @     �D@     �[@      @      @     @P@      *@      L@     �G@     �N@      =@      ,@      @      &@       @      �?      @      5@      @      4@      4@      (@      0@      �?              T@     �m@      @      0@      b@      4@      �@     �C@     �z@     @Z@      @             �F@     �g@      @      "@     �V@      3@     `�@      2@     ps@      L@      @               @     �C@              @      2@             �f@      �?     �T@      $@      @              @      ,@              �?      @              [@      �?      C@       @      @              �?      9@              @      *@              R@             �F@       @                     �B@     �b@      @      @     @R@      3@     �u@      1@     �l@      G@       @              5@      R@       @       @      A@      @      l@      .@      a@      =@                      0@     @S@      �?      @     �C@      *@      ^@       @      W@      1@       @             �A@      I@      �?      @     �J@      �?      V@      5@     �\@     �H@                      :@      E@              @     �@@             @U@      1@     �Z@     �@@                      7@     �D@              @      <@             �M@      ,@      W@      ;@                      @      �?               @      @              :@      @      ,@      @                      "@       @      �?      �?      4@      �?      @      @      "@      0@                              @                      @      �?               @              @                      "@       @      �?      �?      .@              @       @      "@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @1DU�N6@�	           ��@       	                   �5@����թ@f           ,�@                           �?����c�@�           �@                            �?��\��g@�            @v@������������������������       ����(��@?            �]@������������������������       ���e S@�            �m@                          �1@*@��:�@�           ��@������������������������       ��\E.��@q            �g@������������������������       ��»r��@e           �@
                          �7@i��;O)	@�           P�@                           �?���a@�            �u@������������������������       ��	�-(@�             p@������������������������       �s����@8            �V@                           �?���	@�           ��@������������������������       �[��ڃ~@~            �i@������������������������       �)�a�k�	@[           H�@                           @��6|�
@(           ̚@                           �?[;���@�            �y@                            �?��_���@~            �j@������������������������       ��.��n�@            �F@������������������������       ����8@`            �d@                            �?����@}            @i@������������������������       ��J:1�@@            �X@������������������������       ����E�@=            �Y@                           @�����@-           T�@                          �4@(��[F�@�           x�@������������������������       ��(+4�X�?           �|@������������������������       ��3�k�@�            Pt@                            �?���@G           0�@������������������������       ��g���@T            �_@������������������������       �� ���@�            px@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        @     @s@     ��@      >@     �H@     �}@      V@     �@      m@     ��@     0x@      7@      @     �j@      t@      ;@      B@     @t@      Q@     �u@     �g@      x@     0p@      5@      @     �Q@     @c@      &@      1@     `c@      5@     �l@     @U@     �k@      ]@      @              9@     �D@               @      B@       @     @]@      *@     �V@      >@                       @      ,@              �?      "@             �B@       @     �F@       @                      7@      ;@              �?      ;@       @      T@      &@     �F@      6@              @     �F@     @\@      &@      .@     �]@      3@     @\@      R@     �`@     �U@      @              &@      >@       @      �?      .@      �?      C@      6@      B@     �@@              @      A@     �T@      "@      ,@      Z@      2@     �R@      I@      X@     �J@      @       @     �a@     �d@      0@      3@      e@     �G@     @^@      Z@     �d@     �a@      .@             @P@      Q@      �?      @     �H@      @     �E@      5@     �N@      ;@      @              K@     �K@      �?       @     �A@      @      2@      0@     �F@      8@      @              &@      *@              @      ,@      �?      9@      @      0@      @               @     @S@     �X@      .@      ,@      ^@     �D@     �S@     �T@     �Y@      ]@      (@              5@      ;@      �?      @      =@      @      A@      5@     �C@      5@      @       @      L@     �Q@      ,@      "@     �V@     �B@      F@      O@      P@     �W@       @              X@     �j@      @      *@     �b@      4@      �@      F@     0y@      `@       @              9@     �P@      �?             �C@      .@     �a@      @     �U@      @@      �?              *@      ?@                      :@      @      P@       @      F@      :@      �?              �?      @                       @              3@      �?      @      "@                      (@      9@                      8@      @     �F@      �?     �B@      1@      �?              (@     �A@      �?              *@      $@     �S@      @      E@      @                      @      5@      �?              @      �?      D@      �?      3@      @                       @      ,@                      @      "@      C@      @      7@      �?                     �Q@     @b@       @      *@     �[@      @     `@     �B@     �s@      X@      �?             �A@     @T@      �?      @      K@      �?     �u@      0@     �h@      H@                      $@      G@      �?       @      3@             @n@      @     @[@      :@                      9@     �A@              �?     �A@      �?     �Y@      *@     �V@      6@                      B@     @P@      �?      $@     �L@      @     �c@      5@     �]@      H@      �?               @      "@              �?      @      @     �K@      @      ?@      $@                      <@      L@      �?      "@     �I@      �?     �Y@      1@     �U@      C@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @'|d��E@�	           ��@       	                    �?7��R�@�           L�@                           �?z�;
8	@           `�@                            @���Ρ�@�           �@������������������������       ��"x�@           �z@������������������������       �o�˒�@x            �f@                            �?�����	@w           ��@������������������������       �e�r`��	@+           �}@������������������������       ��t$�%{	@L           ��@
                            �?���4c@�           p�@                          �1@�
l�zN@w             h@������������������������       �0q��er @             ?@������������������������       ��ϟ���@f            @d@                           �?�)�gW�@           �x@������������������������       ���(�N�@N            �]@������������������������       �J���@�            `q@                           �?���P�@D           ��@                            �?^�>��Z@p           ��@                           @x��xh��?H            �^@������������������������       �l`��-�?(            �Q@������������������������       �}I�)
@             �J@                          �4@�J<@(           0|@������������������������       ����>O�?�            Pq@������������������������       ����v��@u            �e@                           !@�_�� �@�           ��@                           @q���@�           `�@������������������������       ��m�ȇ�@           `�@������������������������       �g�ӞV�@�            �r@������������������������       �GC7�K@             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        (@     Pr@     h�@      A@     �K@     �z@     �W@     l�@     �m@      �@     �u@      >@      &@     �j@      t@      4@     �E@     0s@     �R@     �x@     �g@     �w@     @m@      ;@      &@      d@     �m@      1@     �B@     �n@     �L@     �m@     �b@     �p@     �f@      8@      @      E@     �V@       @      *@     �W@       @     �_@     �H@     �]@     �K@      @       @      =@     �O@      �?      @     �Q@      @     @T@      C@     @T@      G@      @      �?      *@      <@      �?       @      8@      @      G@      &@      C@      "@               @     �]@     �b@      .@      8@     �b@     �H@     �[@     @Y@     @b@     �_@      2@      @     �N@     �Q@      @      (@     �M@      <@      J@     �N@      O@     �J@      @      @     �L@     �S@      "@      (@      W@      5@     �M@      D@      U@     @R@      &@             �J@     @T@      @      @      O@      2@     �c@      D@     �\@     �J@      @              ,@      @@              @      4@      *@     �F@       @      E@      *@      @                      $@                      �?              (@      �?       @      @                      ,@      6@              @      3@      *@     �@@      @      D@       @      @             �C@     �H@      @      @      E@      @     �[@      @@     @R@      D@                      .@      @                      (@             �J@      @      :@      @                      8@     �F@      @      @      >@      @      M@      =@     �G@      A@              �?      T@     �i@      ,@      (@     �^@      3@     ��@     �H@     @z@      ]@      @              ,@     @R@       @       @      ;@      @      q@      $@     �a@      8@      �?                      0@       @               @      @     �Q@              0@      @                              &@                      �?      @      F@              @      @                              @       @              @       @      :@              $@      �?                      ,@     �L@               @      3@       @     @i@      $@     �_@      2@      �?              $@      @@               @      "@             �a@      @      S@      @      �?              @      9@                      $@       @      O@      @      I@      ,@              �?     �P@     �`@      (@      $@      X@      (@     x@     �C@     `q@      W@       @      �?      O@     @`@      (@      $@     �W@       @     x@     �C@     @q@      W@       @      �?      E@     �X@      @      @     @P@      @     �s@      8@     �h@     �K@       @              4@      ?@      @      @      >@      @     @R@      .@     �S@     �B@                      @       @                      �?      @                       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�chG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @���0@�	           ��@       	                    @�&���@�           ��@                            �?����J�@`           �@                          �<@g�Y���@�           ��@������������������������       �Y�P��@�           ��@������������������������       ���y�� @M            �^@                          �9@�g���@n            �d@������������������������       ��RY�@Q            @^@������������������������       �9lin@             F@
                          �5@W��C�@�           �@                           �?\�U	z3@O           �@������������������������       �k�SP�>@3           �|@������������������������       ��Y8�@           �z@                            �?Nˡ�@=           8�@������������������������       �x�o�2�@[             b@������������������������       ���7���@�            pw@                           �?�ھ3V�@�           ��@                           �?�c	1�@4           �}@                          �9@p�&ᐻ	@�             r@������������������������       ��c�C�7@�            �i@������������������������       �v��.	@3            @T@                          �1@�o��k�@}            �g@������������������������       ��0Z�V @             ?@������������������������       �R��[I@h            �c@                           �?M�S�@�           �@                          �3@�����2@m            `f@������������������������       �� �̋@8             U@������������������������       ���n��3@5            �W@                           @����E|@0           �~@������������������������       ������I@(           �}@������������������������       ��u�B�+@             .@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     X�@     �@@     �K@     �~@      U@     ��@     �g@     h�@     �u@      7@      (@     �i@     �x@      0@      8@      u@     �N@     �@     @`@     ȃ@     `m@      1@      (@     `a@     �f@      &@      1@     �i@      J@      k@      X@     @p@     �b@      ,@      &@     �_@     �d@      &@      1@     `e@      H@     �g@     �V@     �k@      _@      &@      &@      ]@     �c@      &@      .@     �d@      @@     �f@     �R@     �h@     �V@      "@              $@       @               @      @      0@      @      0@      8@     �@@       @      �?      *@      0@                     �@@      @      <@      @     �B@      8@      @              $@      @                      5@      �?      9@      @     �@@      .@      @      �?      @      "@                      (@      @      @              @      "@                     �P@     �j@      @      @     �`@      "@     @~@      A@     Pw@     �U@      @              8@      _@      @      @     �M@      @     �v@      0@     �n@      F@      �?              &@     �L@              @     �C@             @h@      "@     �\@      ?@                      *@     �P@      @              4@      @     `e@      @     �`@      *@      �?              E@      V@       @      �?     @R@      @     �]@      2@     �_@     �E@       @              .@      2@                      .@             �F@      @      :@      4@                      ;@     �Q@       @      �?      M@      @     �R@      *@      Y@      7@       @      "@     �S@     `d@      1@      ?@     �c@      7@     �q@      N@     �j@      \@      @      @      8@     �Q@      (@      "@     �J@      .@     �`@      0@     �U@     �H@      @      @      5@      I@      &@      "@      C@      &@     �J@      *@      D@      @@      @       @      .@      @@      $@      @      =@      @     �J@       @      @@      0@      �?      @      @      2@      �?      @      "@      @              @       @      0@      @              @      4@      �?              .@      @      T@      @     �G@      1@                       @      @                                      0@       @      @       @                      �?      ,@      �?              .@      @      P@      �?      F@      .@              @     �K@     @W@      @      6@      Z@       @     �b@      F@     @_@     �O@       @              ,@      ?@               @      6@              N@      @      B@      "@                       @      $@               @      @              @@              ;@      @                      (@      5@                      1@              <@      @      "@      @              @     �D@      O@      @      4@     �T@       @     @V@     �C@     @V@      K@       @       @      D@      O@      @      4@     �S@       @      V@     �C@     �T@      K@              �?      �?                              @              �?              @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJD~xhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @m�lc�_@�	           ��@       	                    �?G�o��@|           &�@                           �?_��B�@�           x�@                          �3@�"�S'�@7            @������������������������       ���<P��@o            �f@������������������������       �d@ }J6@�            �s@                            �?���-�@o            �c@������������������������       ����x�@$            �K@������������������������       ��{7S&@K             Z@
                            �?t:�ea	@�           �@                           @�
�!sL	@           {@������������������������       ����@|            �g@������������������������       ��uf%�@�            �n@                           @�ƊU�E	@�           L�@������������������������       �:ƃ$	@e           ��@������������������������       ���%�m@U             `@                          �7@�Cy��X@H           ؚ@                          �4@�[�"�@>           ��@                          �1@�`OW��@E           ��@������������������������       �s�n͙�?�             s@������������������������       �)?���@v           �@                           @��yԌ@�            �v@������������������������       �:�(�8@5             T@������������������������       ���e"�-@�            �q@                           @u��,F@
           p{@                           �?�>^�ɶ@�            �q@������������������������       ����L�@A             Z@������������������������       ��aE�e�@n            @f@                          �9@��<��@[            �c@������������������������       �L��ym�@*             R@������������������������       �䜺���@1            @U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �p@     `�@     �C@      J@     p|@      U@     ��@     �k@     H�@     @x@      B@      *@     �g@      u@      =@     �B@     t@     �P@     �w@     �e@     �v@     Pp@      :@             @P@     @X@      @      @     �T@      @     @c@      A@     �a@     �O@      @             �K@     �S@      @      @     �Q@       @     @X@      <@     @Y@     �J@      @               @      ;@              �?      ;@       @     �D@      $@     �F@      4@                     �G@      J@      @      @     �E@              L@      2@      L@     �@@      @              $@      2@              @      *@      �?     �L@      @      D@      $@      �?              �?       @              @      @              3@              0@      �?      �?              "@      $@                      @      �?      C@      @      8@      "@              *@      _@      n@      :@      >@     �m@      P@     @l@     �a@     `k@     �h@      5@      �?     �B@      I@      @      $@     @S@      2@     �Q@     �G@     �O@     �E@      &@      �?      *@      4@              @     �D@      (@      ?@      ,@      5@      :@       @              8@      >@      @      @      B@      @      D@     �@@      E@      1@      "@      (@     �U@     �g@      5@      4@      d@      G@     `c@     @W@     �c@     `c@      $@      @     �Q@      e@      5@      4@     �a@     �D@     �`@     �R@     �b@     `a@       @      @      0@      6@                      3@      @      4@      2@      @      0@       @       @     �S@     @k@      $@      .@     �`@      1@      �@     �H@     z@     �_@      $@             �J@      e@      @      @      T@      @     (�@      8@     @r@     @U@       @             �A@     @\@      @      @      D@       @     @z@      4@      j@     �P@      �?              "@      B@              �?       @              d@       @     @S@      &@      �?              :@     @S@      @      @      @@       @     0p@      2@     �`@      L@                      2@     �K@      @      �?      D@      @      `@      @     �T@      2@      @              @       @       @              �?      @      B@      �?      2@       @      @              .@     �G@       @      �?     �C@      �?     @W@      @     @P@      0@       @       @      :@      I@      @      "@      K@      $@     �V@      9@     @_@      E@       @       @      @      D@              "@      8@      "@     �O@      ,@     �V@      :@                      �?      2@                       @      @      >@       @     �C@      @               @      @      6@              "@      6@       @     �@@      (@     �I@      5@                      5@      $@      @              >@      �?      <@      &@     �A@      0@       @               @      @                      *@              0@      "@      $@       @       @              *@      @      @              1@      �?      (@       @      9@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJPhhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@dj�q�_@�	           ��@       	                    �?X�;��,@m           L�@                           �?Ʌ�a�.@�           ��@                          �3@f��D@�             t@������������������������       �i�G�}�@�             q@������������������������       �@9�'��@              H@                          �1@e�o�ߩ@�            �s@������������������������       ��~:���?X             a@������������������������       ���$��@r            `f@
                           �?���y�]@�           \�@                            �?�^wӴ�@            y@������������������������       �Av�y�~@M             _@������������������������       �_��A;w	@�            @q@                           @.��4��@�           8�@������������������������       ��=�@�            �w@������������������������       �KRF:@�            �x@                           �?|A1lՠ@*           l�@                           �?蚜��@g           ��@                          �<@��
�@�            �p@������������������������       �*롄�@�             k@������������������������       �����{@"            �H@                            �?�	�f�@�            �r@������������������������       �Ɗ��z�@'             Q@������������������������       ��&p6	@�            �l@                            �?t��o�/	@�           �@                           @�q��V	@�           �@������������������������       �����
@4           �}@������������������������       �8%k2�@�            �r@                          �;@�j�iɸ@�           �@������������������������       �����@t           ��@������������������������       ��끭R�	@e            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�       �@@     @r@     �@      ?@      I@      |@      U@     \�@     �m@     x�@     Pt@     �B@      &@      X@     `k@      ,@      0@     `c@      .@     ��@      V@     �x@     @_@      &@             �D@      Q@              @     �C@       @     Pr@      .@      b@      :@      @              ,@      ?@              @      2@       @     �c@      &@     �P@      ,@      @              *@      <@              �?      .@       @     ``@       @      O@      (@                      �?      @              @      @              :@      @      @       @      @              ;@     �B@                      5@              a@      @     �S@      (@                      @      .@                       @             �S@      @      7@       @                      4@      6@                      *@             �L@      �?      L@      $@              &@     �K@     �b@      ,@      (@      ]@      *@     0w@     @R@     �o@     �X@       @      &@      9@     �D@      @       @     �P@      @     @R@      C@     @R@      G@       @              "@      *@                      7@      �?      7@      3@      :@       @       @      &@      0@      <@      @       @      F@      @      I@      3@     �G@      C@      @              >@     �[@      $@      @     �H@      @     �r@     �A@     `f@     �J@                      5@     �L@              @      <@      �?     �b@      .@     �T@      :@                      "@     �J@      $@      �?      5@      @     �b@      4@     @X@      ;@              6@     �h@     `r@      1@      A@     pr@     @Q@     �w@     �b@      z@      i@      :@      �?      K@     �T@               @     �O@      ,@      e@      9@      ]@      A@      @      �?     �@@     �E@               @     �A@             �J@      5@      J@      7@      @      �?      :@     �C@                      <@             �H@      1@      F@      $@      @              @      @               @      @              @      @       @      *@                      5@     �C@                      <@      ,@     �\@      @      P@      &@       @                      @                       @      "@      <@      �?       @      @       @              5@      @@                      4@      @     �U@      @      L@      @              5@     �a@     �j@      1@      @@      m@     �K@     �j@     �^@     �r@     �d@      5@      .@      S@     �]@      @      5@     �W@     �@@     �Y@     �R@     �a@     �T@      @      .@     �H@      S@      @      1@     �P@      <@     �C@     �J@     �P@      K@      @              ;@      E@      �?      @      ;@      @      P@      6@     �R@      =@              @     �P@     �W@      $@      &@     @a@      6@      \@      H@      d@     �T@      2@       @     �E@     @S@      @      @     @\@      *@     �W@      B@      a@     �M@      2@      @      7@      1@      @      @      9@      "@      2@      (@      8@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�
�hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�n9k@�	           ��@       	                    �?�̣Tg�@�           (�@                          �8@��ѐ�@�           Ѓ@                           @
Y �ҍ@B           p�@������������������������       �/�<��@�            �l@������������������������       ���p�L)@�            �r@                          �9@֘�N�@I             [@������������������������       ��O	��@             5@������������������������       ��d�/�C@<            �U@
                           @���l@l           ��@                           �?���:�@�            @v@������������������������       �:��E@�             p@������������������������       �2w�Jt�@4            �X@                          �4@0c�ZӘ @�            �m@������������������������       �ي4#��?Z            `b@������������������������       ���+���@<            @V@                           @l-BVL@�           ��@                          �3@�Ʊ�\	@�           ��@                           @�`!�cS@            �{@������������������������       ��F�Yi@�            �s@������������������������       �5�a��@Y             `@                           @8PKE�~	@�           ��@������������������������       ��=��}~	@�           X�@������������������������       ��iqn�@           �{@                          �7@ Xը|�@�           h�@                           @�a�mw@�           �@������������������������       �"z�@y            �h@������������������������       �����@�           �@                           @ >4��@�            ps@������������������������       ���ɼ�<@K             _@������������������������       ��}��%@j            `g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     0s@     ��@      >@      N@     �{@     �T@     ��@     �l@     8�@     �v@     �@@      �?     @T@     �c@      @      $@      Y@       @     �{@      L@     `q@     �S@      @      �?     �A@     �T@      @       @      K@      @     �o@      @@     �[@     �G@                      =@     �P@      @      @     �E@      @     @m@      5@      W@      :@                      .@      8@      @      @      9@      @     �U@      2@      B@      ,@                      ,@     �E@               @      2@      �?     `b@      @      L@      (@              �?      @      0@              @      &@              5@      &@      2@      5@                       @                      �?      @               @      @      �?      @              �?      @      0@               @       @              3@      @      1@      .@                      G@     @R@       @       @      G@       @     �g@      8@      e@      @@      @             �D@     �C@               @      B@      �?     �U@      1@     �X@      =@      @              =@      B@               @      =@             �L@      *@     �N@      ;@      @              (@      @                      @      �?      =@      @      C@       @       @              @      A@       @              $@      �?     @Z@      @     @Q@      @                      @      ,@                      @             �U@      @     �A@                                      4@       @              @      �?      2@      @      A@      @              1@     @l@     @y@      9@      I@     @u@     �R@     ȁ@     �e@     @     �q@      ;@      *@     `c@     0p@      5@      A@     @m@     �M@      l@     @a@     `k@     @h@      7@      @      A@      M@       @      $@      P@      "@      Z@      E@      Q@      G@      @       @      1@      C@      �?      "@      I@      @     �R@      ;@     �K@     �C@              �?      1@      4@      �?      �?      ,@      @      =@      .@      *@      @      @      $@     @^@      i@      3@      8@     @e@      I@      ^@      X@     �b@     �b@      0@       @      S@      Y@      .@      $@     �\@     �D@     �Q@     �F@     @Y@     �W@      @       @     �F@     @Y@      @      ,@     �K@      "@      I@     �I@      I@     �J@      "@      @     �Q@      b@      @      0@     �Z@      0@     �u@      A@     `q@     �V@      @              J@     �\@      @      &@      N@      ,@     �q@      &@     �h@     �L@       @              2@      A@                      &@      $@      R@      @      ?@      .@       @              A@     @T@      @      &@     �H@      @      j@      @     �d@      E@              @      3@      >@      �?      @      G@       @      P@      7@     @T@      A@       @      @      ,@      @               @      7@              ?@       @      >@      @       @              @      :@      �?      @      7@       @     �@@      .@     �I@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��'KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�|��?@�	           ��@       	                    �?G1��1@           ��@                          �5@vEъ@B           �@                          �3@�k�xe�@�            Pp@������������������������       ��3�H�@w            �g@������������������������       ���xh��@.             R@                            @R�\�L@�            �n@������������������������       �#c���>@j            �e@������������������������       �pϮj؊@3            �R@
                          �5@g f��a@�           `�@                           �?��TD��?E           ��@������������������������       �C�`q��?�            s@������������������������       ��R$t�Z�?�             l@                           @��uRq�@�            @k@������������������������       ��Ɵg}@=            @X@������������������������       �����W�@T            @^@                          �1@�5-�B@�           Ĥ@                           @b0c@�            �v@                           @hP�t3@             H@������������������������       �8%̊]@             ;@������������������������       ���-��?             5@                           @����&�@�            �s@������������������������       �����@�            �q@������������������������       �
�]��@             A@                            @	�=���@�           �@                           @���(jl@�           �@������������������������       ���ʱ	@           �@������������������������       ����`�'@�           �@                           �? R�L<	@�           ��@������������������������       ��5��}�	@�            @n@������������������������       �/0C��i@           |@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     Pr@     ��@     �A@     @Q@     �|@     �S@      �@     �g@     Ј@     �u@      >@      �?     @T@     �f@      @       @     @\@      "@     �}@      A@     �p@     �R@      @      �?      I@      V@      @      @      Q@             �[@      7@     �Z@     �H@      @              ,@     �E@      @              ;@              U@      *@      L@      4@      �?              @     �@@                      8@             �L@      "@      E@      2@                       @      $@      @              @              ;@      @      ,@       @      �?      �?      B@     �F@      �?      @     �D@              :@      $@      I@      =@      @      �?      >@      9@                      <@              5@      @      B@      8@      @              @      4@      �?      @      *@              @      @      ,@      @                      ?@      W@              @     �F@      "@     �v@      &@     `d@      :@                      2@      N@              @      7@      �?     �r@      @     @[@      $@                      $@      @@              @      ,@      �?      f@      @     �M@      @                       @      <@                      "@             �^@      @      I@      @                      *@      @@                      6@       @      Q@      @      K@      0@                      @       @                      &@      @     �C@      @      0@      @                      @      8@                      &@       @      =@       @      C@      "@              *@     �j@     �x@      ?@     �N@     �u@     �Q@      �@     �c@     h�@      q@      9@              .@      J@              @      8@       @     �`@      ,@     �X@      5@                      @      �?                      @              2@      "@      "@      @                      @      �?                      @              @      "@       @      @                                                                      *@              @      �?                      &@     �I@              @      5@       @     �\@      @     @V@      1@                       @      H@              @      ,@             @Z@      @      U@      *@                      @      @                      @       @      $@              @      @              *@     �h@     pu@      ?@     �L@     @t@      Q@     �y@     �a@     �z@     �o@      9@      @      a@     @l@      3@      E@     `l@      G@     ps@     �X@      s@     �e@      (@      @     �T@     �X@      .@      ?@     �`@     �A@     @Y@     �Q@      ]@      Z@      @              K@      `@      @      &@      W@      &@     @j@      <@     �g@     �Q@      @      @      N@     @]@      (@      .@     @X@      6@      Z@      F@     @^@     �S@      *@      @      3@     �C@      &@      @      @@      $@     �C@      @     �A@      A@      @       @     �D@     �S@      �?      $@     @P@      (@     @P@      C@     �U@     �F@      @�t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJbu�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?FNAl�Y@�	           ��@       	                   �<@&B����@            �@                           �?���
@�           ��@                           �?o��%�@�           X�@������������������������       ����n�@�            @h@������������������������       ���;Y!@           �x@                           �?̦ѫj�@Q           �@������������������������       ��JJ%�@�            �m@������������������������       ��b�J>@�            Ps@
                           �?�Zŧ0@5            �T@                            �?DF;�]<@              I@������������������������       ��)���?             &@������������������������       ��ׯ-$�@            �C@                           �?��K�@            �@@������������������������       � ��@�@             1@������������������������       �>��_�@
             0@                            @�ۏa�8@�           �@                           @���僵@�           �@                          �3@�N~�l	@g            �@������������������������       �ݫ��~@�            q@������������������������       ���AѨ	@�           x�@                           @��D:�@t           �@������������������������       ����=5w@�           P�@������������������������       ��Pc@�            �n@                           �?��!� 3	@�           @�@                           �?3����@,             Q@������������������������       ��ϒI@             1@������������������������       ��isP(�@            �I@                           @�8����@�            �@������������������������       ����-
@B            �W@������������������������       ���G�W�@~           (�@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �r@     ��@     �A@      J@     h�@      S@     H�@     �i@      �@      u@      @@             @T@     �e@      @      $@      _@      $@     �z@      A@     �p@     @T@      @             @S@      d@      @      @     �[@       @     0z@      :@     p@      N@      @              B@      R@       @      @     �Q@      @     �o@      0@      Y@      8@      �?              2@      :@       @      @     �A@       @     �G@      $@      C@      (@      �?              2@      G@              @      B@       @     �i@      @      O@      (@                     �D@     @V@      �?              D@      @     �d@      $@     �c@      B@      @              :@      L@                      9@              H@       @      K@      8@       @              .@     �@@      �?              .@      @     @]@       @     �Y@      (@      �?              @      (@              @      *@       @      $@       @      $@      5@                       @      $@              @      "@                      @      @      3@                      �?      @                      �?                               @      �?                      �?      @              @       @                      @       @      2@                       @       @                      @       @      $@      @      @       @                       @      �?                               @      @       @       @       @                              �?                      @              @      @      @                      8@     �j@     @v@      @@      E@     y@     �P@     ��@     �e@     ��@     �o@      <@      *@     �b@     `p@      0@      >@     �p@      D@     �z@     @]@     �y@     `e@      .@      *@     �U@     �`@      ,@      5@     �c@      @@     @a@     �V@     @c@      [@      *@       @      3@     �C@      @      �?      A@      @      Q@      9@     �K@      1@      @      &@      Q@     �W@      $@      4@     �^@      =@     �Q@     @P@     �X@     �V@      @              P@      `@       @      "@     �\@       @     �q@      ;@     p@     �O@       @              F@      Z@               @      S@      @     �m@      4@      f@     �D@       @              4@      8@       @      �?     �C@       @     �H@      @     @T@      6@              &@      P@     �W@      0@      (@     @`@      :@      ]@      L@     @c@      U@      *@      @       @      ,@                      1@      @              ,@      @      @               @      �?       @                              �?              @               @              �?      @      @                      1@      @              &@      @       @               @      L@      T@      0@      (@     @\@      6@      ]@      E@     �b@      T@      *@      @      @      $@      @              .@      @      &@      @      2@      (@      @       @      J@     �Q@      $@      (@     �X@      3@     @Z@      B@     �`@      Q@      "@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJljV8hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?S�[ҫI@�	           ��@       	                    �?&�X�A	@�           ܘ@                          �<@>��\�"@             |@                           �?"���@�            �x@������������������������       �+��lL@w            �f@������������������������       �y뚩�@�            �j@                           �?w�Ѳ�@%             M@������������������������       �-�C�@            �A@������������������������       ��.��)�@             7@
                           �?͹�_��	@�           ԑ@                          �:@(4r1I@            z@������������������������       ���M2��@�            �u@������������������������       ���J��@+            @Q@                           �?2��ρL
@�           ��@������������������������       �oֆ�
@�            �l@������������������������       �~�\�
@8           �~@                           �?�"�2�@�           $�@                          �4@�<_�,�@�           8�@                           @:a6DԺ�?%           �|@������������������������       ������@<            @U@������������������������       ��P%X���?�            �w@                            �?�h7J'`@�            �s@������������������������       ��oN�w@-            @Q@������������������������       ���ށJ@�            `n@                          �5@�%f��@�           ,�@                           @aDp�Z|@I           @�@������������������������       �l�q�@           H�@������������������������       ��GEP@<            �W@                           @0�ps�@�           �@������������������������       ��e�Ǡ@W           ��@������������������������       ��!��"@E            @\@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      t@     ��@      9@      L@      |@     @S@     ��@      k@     8�@     @v@      C@      ,@     `f@     �l@      ,@      >@      n@     �I@     �j@      a@     �o@     �h@      ?@              J@     �R@               @      O@       @     �U@      9@      V@     �G@      @              I@      O@              @     �H@       @      U@      5@      U@      =@      @              7@      @@              @      3@       @      E@      (@      >@      *@      @              ;@      >@              �?      >@              E@      "@      K@      0@      @               @      (@              @      *@               @      @      @      2@                              &@               @      @              �?      @      @      (@                       @      �?              �?      $@              �?      �?      �?      @              ,@     �_@     `c@      ,@      6@     @f@     �H@      `@     �[@     �d@     �b@      9@      �?      B@     �M@       @      @      R@       @      Q@     �B@     �N@     @P@       @             �@@     �K@       @      @      O@      @     �N@      =@      J@      E@       @      �?      @      @              �?      $@      @      @       @      "@      7@              *@     �V@      X@      (@      .@     �Z@     �D@     �N@     �R@     �Z@     @U@      7@       @      6@      E@      @      @      >@      4@      5@      5@      7@      A@      @      &@     @Q@      K@       @      "@      S@      5@      D@     �J@     �T@     �I@      1@       @     �a@     0s@      &@      :@     @j@      :@      �@     @T@     @�@     �c@      @              A@      U@       @      @     �E@      "@     �v@       @      i@      :@      @              4@     �C@              @      6@             `n@      @     @]@      (@       @              "@      @              �?      @              <@      �?      <@      @                      &@      A@              @      .@             �j@       @     @V@      @       @              ,@     �F@       @              5@      "@     �]@      @     �T@      ,@      �?                      @       @               @       @      =@              4@      �?      �?              ,@     �C@                      *@      @     @V@      @     �O@      *@               @     �Z@     �k@      "@      5@     �d@      1@     p{@     @R@      v@     �`@      @             �C@     ``@      @      &@     @R@      $@     0s@      :@     �m@     �O@      @             �@@     �]@      @      @     �P@       @     �q@      7@     �k@      G@      �?              @      *@              @      @       @      9@      @      0@      1@       @       @      Q@      W@      @      $@     �W@      @     �`@     �G@      ]@     �Q@      �?       @     �G@     �R@      �?      $@      S@      @     �\@      >@     �Y@     �P@                      5@      2@      @              2@      �?      1@      1@      ,@      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ'Yw<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@>G��Zi@�	           ��@       	                   �1@)�����@U           ��@                           �?�}l�:z@m           8�@                            �?�+U��@i            �c@������������������������       �01���@5            �T@������������������������       �t��;�@4            �R@                            �?{����.@           �x@������������������������       ���7=zV @�             l@������������������������       ��N� @s            @e@
                            @�'��@�           `�@                           �?�H�(Y�@�           ��@������������������������       ��ڹ�Ȣ@J           ��@������������������������       �r�`G��@�           ��@                           �?�<�wd�@           �z@������������������������       �N����M@P            �`@������������������������       �(��4�p@�            pr@                          �:@��]S�@K           (�@                           �?Ή�ی8@�           <�@                          �7@�f�L�	@W           �@������������������������       �=�G�N@�            �m@������������������������       �*v��2�@�            `s@                           @�b�c}@�           `�@������������������������       �����@R           �@������������������������       ���#�@5            �R@                           �?J_�f*	@m           ؁@                           �? ���	@�            t@������������������������       ��6�-P@G            �]@������������������������       �?��*�	@�            @i@                           @p�g=�@�            @o@������������������������       �$,�2E@G            �]@������������������������       �bb���@U            ``@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     �@      @@     �L@     �|@     �R@     ��@     �m@     x�@     �u@      A@       @     �_@     �r@      .@      4@     �j@      A@     @�@     �X@     @@      e@      (@      �?      :@     @R@      �?      @      D@       @     �l@      1@     �]@      C@      �?      �?      &@      8@      �?              8@       @      C@       @      9@      7@              �?      @      2@                      &@       @      .@      �?      1@      *@                      @      @      �?              *@              7@      @       @      $@                      .@     �H@              @      0@             �g@      "@     �W@      .@      �?                      :@              @      $@              ]@      @     �G@      *@                      .@      7@                      @             �R@       @     �G@       @      �?      @     @Y@      l@      ,@      .@     �e@      @@     @|@     �T@     �w@     ``@      &@             �T@     �d@      "@      @     �^@      1@      v@      P@     `q@     �V@      @             �A@     �P@      @      �?      M@      @     @g@      C@     �W@      C@      @             �G@     �X@      @      @      P@      $@      e@      :@      g@      J@       @      @      3@      M@      @      "@      J@      .@     �X@      2@     �Y@     �D@      @              &@      .@              @      $@              I@      @      <@      ,@              @       @     �E@      @      @      E@      .@      H@      .@     �R@      ;@      @      &@     �e@     @o@      1@     �B@     �n@     �D@     �r@     @a@     �s@     �f@      6@      @     @\@     �g@      &@      8@     �c@      8@     `m@     �R@      k@     @Y@      1@       @     �P@     @^@       @      1@      T@      &@     �Q@      H@      Q@     �D@      .@       @     �A@     �J@      �?      @     �A@      @      5@      *@     �B@      9@      @              ?@      Q@      @      &@     �F@       @     �H@     �A@      ?@      0@      "@       @     �G@     �Q@      @      @     @S@      *@     �d@      :@     �b@      N@       @       @      B@      O@      �?      @     @Q@      $@     @c@      (@      a@      L@                      &@       @       @               @      @      &@      ,@      &@      @       @      @      O@     �M@      @      *@     �V@      1@      Q@      P@     �X@     @T@      @      @      D@     �A@      @       @     �F@      *@      A@     �A@      E@      K@      @       @      @      $@               @      2@       @      5@      &@      8@      3@      @      @      A@      9@      @      @      ;@      &@      *@      8@      2@     �A@      �?              6@      8@      @      @     �F@      @      A@      =@     �L@      ;@                      @      *@      @      @      0@       @      1@      7@      6@      ,@                      1@      &@              �?      =@       @      1@      @     �A@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��;ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��=k�Y@�	           ��@       	                   �2@_�`���@W           ֠@                           �?��U!Ea@&           �|@                           @���!r@p             d@������������������������       ��`��@S             _@������������������������       � 6��@             B@                            �?���<��@�            �r@������������������������       �ޠ!�Zq@=             X@������������������������       �6��B�@y            @i@
                          �;@�U�l	@1           ��@                           �?f�xj%	@_           \�@������������������������       ��?��@�            �x@������������������������       ��I��	@b           p�@                           �?"��n��	@�            �t@������������������������       �:�Θq�@A            �Z@������������������������       �% ���	@�             l@                          �3@i�(T4@L           x�@                           @S��M.@�           ��@                          �2@B�>��7 @X           8�@������������������������       ����:�?�            �y@������������������������       �ҙA�X@a            �a@                            �?�sV�P�@y             i@������������������������       �0m��}�?            �K@������������������������       �Y('�Uv@Z            @b@                           @2�%e��@{           p�@                           @4�	h1@�           Ȅ@������������������������       ��ꪎ@           �z@������������������������       �m��@�            �m@                           �?v��J|�@�            Pu@������������������������       �Bs��A@b            �b@������������������������       �I1�H@y            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@      r@     `�@      A@      N@     pz@      S@     �@      k@     ��@      x@      <@      8@     �h@     �u@      <@      D@     �q@      L@     0w@      f@      v@     �p@      3@       @      =@     �R@              �?     �G@       @     �a@      ;@     �V@      F@      �?       @       @      ?@                      4@      �?      K@      (@      1@      ,@      �?              @      7@                      2@             �F@      "@      ,@      "@               @       @       @                       @      �?      "@      @      @      @      �?              5@     �E@              �?      ;@      �?     �U@      .@     �R@      >@                      @      2@                      @      �?      >@      @      4@      (@                      .@      9@              �?      7@              L@      $@      K@      2@              6@     �d@     �p@      <@     �C@     �m@      K@     �l@     �b@     Pp@     �k@      2@      (@     �`@     �l@      7@      ;@      i@      D@      j@     @]@     `k@     �a@      *@             �F@     �P@       @      @      ?@       @     �W@      2@     �V@     �C@      �?      (@     �U@     �d@      5@      8@     @e@      C@     �\@     �X@      `@      Z@      (@      $@     �A@     �C@      @      (@     �B@      ,@      6@      @@      E@     @S@      @      @      $@      *@              @      0@              @      &@      .@      6@       @      @      9@      :@      @      @      5@      ,@      0@      5@      ;@     �K@      @      �?      W@     �j@      @      4@     @a@      4@     P�@     �D@     �{@     �^@      "@              :@     �V@              "@     �D@      �?     `v@       @      g@      @@       @              2@     �R@                      9@      �?     �p@      @      a@      9@                      (@      L@                      $@      �?      k@      �?     �W@      2@                      @      2@                      .@              J@      @     �D@      @                       @      1@              "@      0@             �V@      @      H@      @       @                      @                      �?             �@@              0@                               @      (@              "@      .@             �L@      @      @@      @       @      �?     �P@     @^@      @      &@     @X@      3@     @r@     �@@     pp@     �V@      @      �?      H@     �R@              �?      M@      @      l@      0@     �f@      J@      @      �?      B@     �D@              �?     �F@      @      `@      $@     �\@     �C@      @              (@     �@@                      *@             �W@      @     �P@      *@                      2@     �G@      @      $@     �C@      ,@      Q@      1@     �T@      C@       @               @      6@       @       @      2@      @      ;@       @      ?@      3@                      $@      9@      @       @      5@      @     �D@      "@     �I@      3@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJs��yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?,��?h@�	           ��@       	                    �?�N$��Z	@�           �@                           �?���b:@/           �|@                           �?�~!���@s            �d@������������������������       �#�6�}�@4             S@������������������������       ��ArH��@?             V@                            �?{#u��@�            �r@������������������������       �\��-T@`            `b@������������������������       ��a@�@\             c@
                           �?�[\yt�	@�           ��@                            �?�����$@           py@������������������������       �Qq�:�@I            �\@������������������������       �#1�O@�            @r@                           @@ ���8
@�           ��@������������������������       ���%�
@�            �@������������������������       �_��˂@	             4@                          �5@��3_�*@�           �@                           @z)~aMm@o           ȕ@                           @���+i�@w           P�@������������������������       ���z�{@�            �w@������������������������       �)�˿f@�            �i@                           �?�Q��~@�           @�@������������������������       �����Α�?�            �q@������������������������       �%M_R��@@           P�@                           @��o6�@?           �@                          �=@�w�m@�           ��@������������������������       �0�	�@t           ��@������������������������       �z['Vb@0            @R@                           �?��L���@�            �o@������������������������       �HR�|�b@K            @_@������������������������       ���#�K(@P             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �q@     @�@      ?@      K@     |@     �T@     h�@      o@     ��@     v@      =@      7@     `d@      m@      5@      @@     �n@      G@     �l@     @b@     �n@     `g@      5@       @     �D@      P@      �?      $@     �K@      @     @[@      :@     @X@      I@      @       @      &@      5@                      5@              H@      @      E@      ,@      �?       @      @       @                      ,@              9@      @      .@      @                      @      *@                      @              7@      �?      ;@      $@      �?              >@     �E@      �?      $@      A@      @     �N@      6@     �K@      B@       @              ,@      0@      �?      @      0@              9@      $@      A@      9@       @              0@      ;@              @      2@      @      B@      (@      5@      &@              5@     �^@      e@      4@      6@     �g@     �D@     �^@      ^@     �b@      a@      2@       @      <@      R@      @      &@     �R@      @      O@     �B@      L@     �J@      �?              @      0@              @      <@       @      3@      4@      ,@       @               @      9@      L@      @      @     �G@      @     �E@      1@      E@     �F@      �?      3@     �W@     @X@      .@      &@     �\@      B@      N@     �T@     �W@      U@      1@      (@     @W@     �W@      .@      &@      \@      B@      N@      T@     �W@     �T@      .@      @      �?      @                       @                      @               @       @      �?      _@     �s@      $@      6@     �i@      B@     0�@     �Y@     8�@     �d@       @             �J@     @g@      @      $@     �\@      &@     P�@      F@     Pu@     �Q@      @              9@     �W@               @      I@      &@     �j@      ?@      ]@     �E@       @              4@      F@               @     �@@       @     `d@      (@     �R@      7@                      @      I@                      1@      @     �H@      3@      E@      4@       @              <@      W@      @       @     @P@             `u@      *@      l@      ;@      @              (@      ;@              @      (@             �c@      @     @P@       @      @              0@     @P@      @      @     �J@             @g@      @      d@      9@      �?      �?     �Q@     �`@      @      (@     �V@      9@     �k@     �M@     @j@      X@       @      �?     �L@     �V@      �?       @     �P@      *@     �f@      C@      c@      N@       @      �?      G@     @T@      �?      @     �H@      &@     `e@      ;@     �b@     �K@      �?              &@      $@              �?      1@       @      &@      &@      @      @      �?              ,@      E@      @      @      8@      (@      C@      5@      M@      B@                      @      ;@       @       @      &@      @      1@       @      =@      1@                       @      .@      @       @      *@      @      5@      *@      =@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�����K@�	           ��@       	                     @W�)4�@           ��@                            �?��$W@H           x�@                            �?���K�@�           ��@������������������������       ��.��c}@�            �u@������������������������       ��$s��@�            @w@                          �3@��8w@�            �k@������������������������       ��.��0 @7            �W@������������������������       �-@�ș�@P            �_@
                           �?R��~jV@�            �t@                           �?,x�@w            @h@������������������������       �f�/1:�@            �E@������������������������       ��y�]w�@Z            �b@                           @�R�Ǌ�?Z            �a@������������������������       ��ϷW���?+            �Q@������������������������       ���$ȱ�?/            @Q@                          �3@*(�K0@�           ��@                           @\PK��@;           ��@                          �1@�ǀ
5�@-           �@������������������������       �H�NiZ@�            t@������������������������       �t�ȃ�@]            �@                             @��P}�@             5@������������������������       ��t�I�|�?             "@������������������������       ��D=�U�@             (@                          �9@���R��@�           X�@                           @�_"s�j@           В@������������������������       �r��8@�           �@������������������������       �a�AS�@             G@                            @'@��Pf	@t           �@������������������������       �VƂ��@�            `u@������������������������       �#�1���	@�            �i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     X�@      @@     �P@      z@     �V@     `�@     �j@     H�@      v@      <@             �V@     �d@       @      (@     �W@      .@     0|@      D@     �s@     @T@      @              O@     �]@      @      @     �P@      ,@     �u@      <@     �m@     �J@      @             �H@      X@      @      @     �J@      &@     @o@      4@     �f@     �F@      @              6@      I@      @       @      6@      @     �_@      @     �U@      9@      @              ;@      G@      @      @      ?@      @      _@      ,@     @X@      4@       @              *@      6@                      ,@      @     �X@       @     �J@       @      �?              �?      @                      @      �?     �J@      @      2@      @      �?              (@      2@                      $@       @     �F@      �?     �A@      @                      <@      H@       @      @      ;@      �?     �Y@      (@     �S@      <@                      ;@     �C@       @      @      5@      �?      C@      $@      @@      3@                       @      (@                       @              .@      �?      $@      �?                      9@      ;@       @      @      3@      �?      7@      "@      6@      2@                      �?      "@               @      @             @P@       @      G@      "@                      �?      @                      @              <@              9@      @                               @               @      @             �B@       @      5@       @              ,@     �i@     Px@      8@     �K@     @t@     �R@     H�@     �e@     x�@     �p@      6@      @      D@     �a@      �?      ,@     @U@      &@     @p@     �K@      i@     @R@       @      @      D@     @a@      �?      ,@     �T@      $@      p@     �K@     @h@     @Q@      �?      �?      *@     �F@              @      6@             �^@      2@     @T@      0@               @      ;@     @W@      �?      &@      N@      $@      a@     �B@     @\@     �J@      �?       @               @                      @      �?       @              @      @      �?                                                               @              @      @               @               @                      @      �?                      @              �?      "@     �d@      o@      7@     �D@     �m@      P@     Pr@      ^@     pt@     �h@      4@      @     �Z@     �h@      &@      @@     @f@      D@     �k@     @P@      m@     @Z@      *@      @     @X@      h@      "@      @@     �e@     �B@     �j@      L@     �l@      Y@      *@      �?      $@      @       @              @      @      @      "@      @      @              @      N@     �J@      (@      "@     �N@      8@     @R@     �K@     �W@     @W@      @       @      @@      C@      @      @      F@      *@      D@      ?@     @Q@      N@      @       @      <@      .@      @      @      1@      &@     �@@      8@      :@     �@@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ6�?hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@��h:@�	           ��@       	                    @.��_@@_           ��@                            �?�9e��0@�           t�@                           �?�n�f@           `|@������������������������       �0��ʨ2@�             t@������������������������       ���	�av@Y            �`@                           �?>W$m@�           \�@������������������������       �I�4��@�           @�@������������������������       �u{&^\N@�            �t@
                           �?T�$c��@�           ��@                          �4@�Mx�@�           @�@������������������������       �v����7@.           �}@������������������������       ���n+�@�            �p@                          �7@|�>�c@�           ��@������������������������       �*�s�@�           `�@������������������������       ��n	 @             H@                           �?�q$�8	@A           @�@                           �?�{�7�	@8           0@                          �<@��mO�@Y            �b@������������������������       �[�ۻǸ@6            @T@������������������������       �O~cn/@#             Q@                           �?��0A�
@�            �u@������������������������       ����F�	@N             ^@������������������������       � �;{	@�            �l@                            @�� �X@	           Py@                            �?��T!�@�            @s@������������������������       �	ʾ�P�@;            @U@������������������������       ��Җ@�            �k@                           �?����W@9            @X@������������������������       �罨, o�?             B@������������������������       ����!�e@'            �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �s@     x�@      :@      E@      }@      U@     H�@      j@     h�@     �u@      <@      "@     @k@     �}@      2@     �@@     �u@      H@     �@     �\@     ��@      l@      0@      "@     �c@     p@      *@      =@     �l@      A@     �r@     �X@     pq@      b@      ,@             �E@      R@              @     @P@      "@     @Z@     �A@     �U@      :@       @              C@     �H@              @      I@      @     �N@      ?@      O@      1@      @              @      7@                      .@      @      F@      @      9@      "@      @      "@     �\@      g@      *@      9@     �d@      9@     @h@     �O@      h@     �]@      @      "@     �U@     �^@      $@      4@     @`@      4@     �\@      F@     �\@      Y@      @              =@      O@      @      @      B@      @      T@      3@     �S@      2@                      N@     �k@      @      @      ]@      ,@     ��@      0@     �v@     @T@       @             �@@      \@       @      @     @T@      "@      q@      @     �f@      F@       @              5@      Q@       @      @     �@@             @i@      @     �\@      =@                      (@      F@                      H@      "@     �Q@      �?     @P@      .@       @              ;@      [@      @      �?     �A@      @     `r@      $@     �f@     �B@                      9@      [@      @      �?      <@      @      q@       @     �d@     �A@                       @                              @              6@       @      *@       @              *@      X@     �\@       @      "@     �]@      B@      a@     �W@     �a@     @_@      (@      *@     �K@     �P@      @       @     �O@      =@     �G@     @P@      N@     �T@      &@      �?      7@      5@                      >@       @      *@      (@      ;@      3@      �?      �?      *@       @                      *@       @      (@       @      5@       @      �?              $@      *@                      1@              �?      @      @      1@              (@      @@     �F@      @       @     �@@      ;@      A@     �J@     �@@     �O@      $@       @      @      6@      @       @      $@      (@      @      2@      &@      6@      @      @      <@      7@      @              7@      .@      =@     �A@      6@     �D@      @             �D@      H@       @      @      L@      @     @V@      =@     �T@     �E@      �?             �@@     �E@      �?      @      I@      @      G@      5@     �P@     �@@      �?              @      &@                      *@              ,@      @      8@      $@      �?              <@      @@      �?      @     �B@      @      @@      ,@      E@      7@                       @      @      �?              @             �E@       @      0@      $@                                                                      6@      @      "@       @                       @      @      �?              @              5@      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��oYhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?|38�zF@�	           ��@       	                    �?��T:*I	@�           h�@                           �?�q��x@s           ��@                          �6@�C�J�a@r            �d@������������������������       ��Z���@G             Z@������������������������       �����r/@+            �N@                           @s]����@           �x@������������������������       �皵`,�@�            @v@������������������������       �JS���@            �E@
                           �?<�P$B�	@r           0�@                            �?�/vG�	@�            pw@������������������������       ��:���~	@u            �h@������������������������       ��F.�#�@s            `f@                            @��*g�J	@�           x�@������������������������       �����%l	@�            �s@������������������������       ���_�4�@�            ps@                           �?�2r\��@�           ^�@                           @Y�����@�           ؇@                            �?��1�	�@l             d@������������������������       ��`�զ @+             O@������������������������       ��#��@A            �X@                           �?m��q� @r           ؂@������������������������       ��d�E @�            �t@������������������������       �tT`;�@�             q@                           @��|	@�           И@                           �?��^�@�            px@������������������������       �$��@[ @             5@������������������������       �Ț�sPm@�             w@                           @S�y��/@�           ��@������������������������       �`ַ8�@�           <�@������������������������       ����PB@             >@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     ��@      :@      H@     p|@      V@     ȏ@     �j@     ��@     0u@     �@@      2@     �e@     �m@      5@      :@     p@     �H@      k@     �`@     �k@     �f@      8@              I@     @Y@      �?      &@      Z@      @     @\@     �@@     @S@     �M@       @              4@      ;@                      7@             �G@      @     �A@       @                      @      5@                       @             �B@      @      :@      @                      0@      @                      .@              $@      �?      "@      @                      >@     �R@      �?      &@     @T@      @     �P@      <@      E@     �I@       @              7@      Q@      �?      $@     �Q@      @      P@      8@     �D@     �F@      @              @      @              �?      &@               @      @      �?      @      @      2@     �^@      a@      4@      .@      c@      E@      Z@     @Y@     @b@      _@      0@      @     �G@      Q@      *@      @     �E@      6@      ;@      A@      B@     �P@      "@       @      8@     �@@      @       @      1@      $@      4@      ;@      "@     �C@      @      @      7@     �A@      @      �?      :@      (@      @      @      ;@      <@       @      (@     �R@     @Q@      @      (@     �[@      4@     @S@     �P@     �[@     �L@      @      @     �E@      A@      @      &@     �M@      "@      >@      ;@     �J@     �@@      @      @      @@     �A@       @      �?     �I@      &@     �G@      D@     �L@      8@      @             �a@     `v@      @      6@     �h@     �C@      �@     �S@     ��@     �c@      "@              :@     �Y@              @     �D@       @     �u@      0@     `g@      A@                      "@      0@               @      0@       @      L@      @     �G@      @                              &@               @      @      �?      6@              4@                              "@      @                      $@      �?      A@      @      ;@      @                      1@     �U@              �?      9@      @      r@      &@     �a@      ;@                      @      H@              �?      (@       @     �e@      @      O@      1@                      $@      C@                      *@      @      ]@      @     �S@      $@                     @]@      p@      @      3@     �c@      ?@     `|@      O@     @v@     �^@      "@             �B@      U@       @      "@      I@       @     �R@      @@      P@      =@       @               @      @              @      @                                      �?                     �A@     @S@       @      @     �E@       @     �R@      @@      P@      <@       @              T@     �e@      @      $@     �Z@      7@     �w@      >@     @r@     @W@      @             @R@     @e@       @      $@     �Y@      *@     �w@      ;@     0r@      W@      @              @       @      �?              @      $@              @      �?      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��MhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�NmQ�x@�	           ��@       	                    �?�Q�)+	@	            �@                           @*BNK@�           Ђ@                            �?Y�+�[@�            �x@������������������������       ��=�Q@�             l@������������������������       �G�k@j             e@                          �9@_۪��@�             j@������������������������       �g5.A@g            �b@������������������������       ��1M���@&            �M@
                          �;@<O�I��	@}           0�@                           @��W��9	@            �@������������������������       ���sz�@�           ��@������������������������       �/��H�%	@y            �h@                           @�<���$
@z            @h@������������������������       �^,�?�	@m            �e@������������������������       ���ю@             5@                          �5@��To@�           �@                          �1@#�qS�@�           ��@                           @��bL��@           `|@������������������������       ���c�cc@
            {@������������������������       ���Ss* @             6@                          �4@��l��@t           P�@������������������������       �t�f���@�           ��@������������������������       ��eA��H@�            �n@                           @T<.�S7@(           Ȋ@                           @��<�q�@�           �@������������������������       ��e�!wR@�            0v@������������������������       �\k��\@�            �q@                          �>@�M��'�@�             k@������������������������       ��1��v5@�            �h@������������������������       ��~�.�@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     q@     @�@     �C@     �L@     �|@     �S@     P�@     �j@     H�@      y@     �@@      5@     �b@     �n@      3@      @@      l@     �@@      m@      b@     @o@      l@      :@      @      D@     @Z@       @      "@     @T@      "@      `@     �B@      [@     �S@       @      @      5@     �P@      �?      �?      J@      @     �X@      5@      T@      F@       @       @      (@      A@                      9@      @      I@      ,@      J@     �@@              �?      "@      @@      �?      �?      ;@      �?      H@      @      <@      &@       @              3@     �C@      �?       @      =@      @      >@      0@      <@      A@                      2@      >@      �?      @      7@      @      9@      $@      0@      1@                      �?      "@               @      @      �?      @      @      (@      1@              2@      [@     �a@      1@      7@     �a@      8@     @Z@     �Z@     �a@     @b@      8@      @      V@     @[@      .@      .@     �_@      *@      X@     �W@     @^@     �Y@      2@      @     �R@     �R@      "@      (@      X@      $@     �R@      L@     �Y@     �U@       @      �?      *@     �A@      @      @      ?@      @      6@     �C@      2@      1@      $@      ,@      4@      @@       @       @      0@      &@      "@      (@      5@     �E@      @      @      3@      =@       @       @      ,@      &@      @      &@      4@      E@      @      @      �?      @                       @              @      �?      �?      �?      �?       @     @_@      s@      4@      9@     �m@      G@     �@     �Q@     x�@     @f@      @             @Q@     `g@       @      0@     �]@      2@     Ё@      B@     `u@     �U@      @              0@     �J@              @      :@              i@       @      ^@      7@      �?              0@      J@              @      :@             @h@       @      ]@      .@      �?                      �?               @                      @              @       @                     �J@     �`@       @      $@      W@      2@     w@      <@     �k@      P@      @              H@     �U@       @      @     �Q@      (@     �q@      8@     �d@     �J@                      @      H@              @      6@      @     �T@      @      M@      &@      @       @      L@     �]@      (@      "@      ^@      <@     �h@      A@      g@     �V@       @       @      H@     �U@              @     �U@      7@     @e@      8@     �`@      O@       @       @      .@      D@               @     �G@      0@     �\@      @     @R@     �C@                     �@@     �G@               @      D@      @     �K@      2@     �M@      7@       @               @      @@      (@      @     �@@      @      =@      $@     �J@      =@                      @      ?@      @      @      @@      @      =@      "@      J@      7@                      �?      �?      @              �?      �?              �?      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@�UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�҇�2@�	           ��@       	                    �?���:@T           ��@                           @���H�@�           ��@                            �?s;Y���@�            Pv@������������������������       �I�Y��@M             ^@������������������������       ��m�/�7@�            �m@                          �0@F߶��]�?           py@������������������������       �V��?            �H@������������������������       ��?��L��?�            `v@
                           �?��p�ge@c           ��@                           @ 8��>�@H           �@������������������������       �-�A��@�            �t@������������������������       ��M���	@j            �f@                            �?��W�@            �@������������������������       �P*᧕�@�             l@������������������������       �,��;�@�            �@                           �?t*ط��@B           ��@                           �?�)Ux�@+           `~@                           �?�!�P�@�            �n@������������������������       ���>�B@4            @U@������������������������       ��p���@`            �c@                          �>@���~3@�            @n@������������������������       �<v��O�@�            @l@������������������������       �+�%W�@
             0@                          �8@�%tA	@           �@                           @�����G@l           P�@������������������������       ��<S�8	@�            �v@������������������������       �0L�}3M@�            �k@                           @fǷ���	@�           ؅@������������������������       �iJ��_1
@           �|@������������������������       ���zB$�@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �t@     ��@      8@     �L@     �{@     �Q@     h�@     `l@     0�@     �u@      8@      (@      a@     �s@       @      3@      g@      8@     �@      U@     �|@     @b@      @             �E@     �X@      �?      @     �G@      @     u@      4@     �e@      @@      �?              =@      H@      �?      @      =@       @     �\@      1@     @W@      4@      �?              @      7@                      @      �?     �@@      @      E@      @                      :@      9@      �?      @      7@      �?     @T@      (@     �I@      *@      �?              ,@     �I@               @      2@       @     �k@      @     �T@      (@                              .@                      �?              3@              $@      @                      ,@      B@               @      1@       @     �i@      @      R@       @              (@     @W@     �k@      @      ,@     @a@      4@      y@      P@      r@     �\@      @      (@      K@      Q@       @      "@     �S@      (@     �R@     �C@     �X@     �N@      @      @      ?@      E@       @      @      L@      @      E@      7@     @S@      E@              @      7@      :@              @      6@      @     �@@      0@      5@      3@      @             �C@      c@      @      @      N@       @     pt@      9@     �g@     �J@                      &@      =@               @      4@      �?     �Y@      @      A@      3@                      <@     �^@      @      @      D@      @      l@      4@     �c@      A@              &@     �h@     �k@      0@      C@     �o@      G@     ps@     �a@     ps@     �i@      1@              H@     @Q@      �?       @      I@      $@     �[@     �@@     @]@     �F@      �?              A@     �C@      �?       @      A@      �?      @@      3@      I@      ?@      �?              5@      @                      *@              4@       @      1@      @                      *@      @@      �?       @      5@      �?      (@      1@     �@@      :@      �?              ,@      >@                      0@      "@     �S@      ,@     �P@      ,@                      &@      =@                      ,@       @      S@      "@     �P@      (@                      @      �?                       @      �?       @      @               @              &@     �b@     @c@      .@      B@     �i@      B@      i@     �[@     @h@     �c@      0@      @     �P@     �S@      @      $@      X@      0@     �]@      ?@     �X@      L@      @      @     �I@      H@      @      "@     @Q@      (@     �H@      9@      J@      B@      @              0@      >@      �?      �?      ;@      @     �Q@      @      G@      4@               @     @T@      S@       @      :@     @[@      4@     �T@     �S@      X@     �Y@      &@       @      N@     �I@      @      4@      Q@      2@     �F@     �P@     �C@     �P@      &@              5@      9@       @      @     �D@       @     �B@      (@     �L@      B@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJkk-OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@.��9Z@�	           ��@       	                    �?ť�vJK@t           4�@                           @oN9U@�           ��@                           �?�Z�B@�             q@������������������������       �N�)�b�@R            �^@������������������������       ��hk}@b            �b@                           @�}c�ҿ�?�            `v@������������������������       ����Gk�?�            `n@������������������������       �v҅���@H            �\@
                           @	��;su@�           T�@                           �?}�-�@�           ��@������������������������       ���;��@�            �y@������������������������       ��O��]@�            �u@                           �?2_odEs@            z@������������������������       � Cv�F@�            @i@������������������������       ���ܑZ@�            �j@                           @еO�X�@;           x�@                          �<@�1�4@�           ��@                           �?����@�           �@������������������������       �8���@)           �|@������������������������       ���cNa@�           ԑ@                           @����`	@�            Pr@������������������������       �3��o�T	@�            �j@������������������������       ���4�;@2             T@                          �:@�,�L�	@�            `j@                           @d��"\�@b            �a@������������������������       ���L��@<            �T@������������������������       ���}*�@&             M@                            @�=���@-            �Q@������������������������       �j�<��X@$            �J@������������������������       ������=@	             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      r@     H�@      =@      P@     �z@     �Y@     ��@     @l@     �@     �v@      5@      @     �T@     @n@       @      6@      d@      8@     ��@     @X@      x@      b@      @              6@     �U@              "@      C@      @     �q@      1@     `b@      <@      �?              0@      C@              @      8@      @      T@      .@      R@      5@                      @      3@              @      2@      @      D@      (@      0@      @                      &@      3@               @      @              D@      @      L@      ,@                      @      H@              @      ,@              i@       @     �R@      @      �?              @      A@                       @             �b@             �G@                              �?      ,@              @      @              J@       @      <@      @      �?      @     �N@     �c@       @      *@     �^@      5@     �u@      T@     �m@     @]@      @      @      I@     �[@       @       @     @X@      5@     `d@     �R@      `@     �V@      @      @      B@     �E@      @      @      N@      0@     @Q@     �D@     @P@     �P@      @              ,@     �P@       @      @     �B@      @     �W@     �@@      P@      8@                      &@      G@              @      9@             @g@      @     �[@      ;@                      @      2@              @      .@             �W@       @      I@      0@                       @      <@              �?      $@              W@      @      N@      &@              *@     �i@     ps@      5@      E@     �p@     �S@     �w@      `@     z@     �k@      1@      @     �e@     pq@      3@      E@     �m@      Q@      v@      Z@      y@     �i@      &@      @     @b@     `n@      ,@      =@     �h@      K@      t@      T@     pv@     @b@      "@             �C@     �S@      @      @      I@      (@      ^@      "@     �\@     �@@              @     �Z@     �d@      &@      9@     �b@      E@     @i@     �Q@     �n@     @\@      "@      �?      =@      B@      @      *@      D@      ,@      >@      8@     �D@      M@       @      �?      9@      8@      @      (@      :@      *@      $@      8@      6@      I@       @              @      (@      �?      �?      ,@      �?      4@              3@       @               @      >@      @@       @             �@@      $@      >@      9@      1@      2@      @      �?      8@      =@       @              .@      "@      9@      &@      $@       @      @      �?      *@      8@                      *@       @      $@       @      @      @      @              &@      @       @               @      @      .@      @      @      @       @      @      @      @                      2@      �?      @      ,@      @      $@              �?       @       @                      .@      �?      �?      ,@      @      $@              @      @      �?                      @              @                                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ{Ǽ6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�-×�7@�	           ��@       	                    @y����K@e           �@                           �?S�@�           �@                           �?�|=��@�            w@������������������������       ����@h            @e@������������������������       ��w�\W@|            �h@                           �?��h��@�           ��@������������������������       ��h4[�N@6           @~@������������������������       �f	Hʪ�@�            �m@
                          �3@����8t@�           �@                           @�0�q2@�           X�@������������������������       �M�&s���?�             w@������������������������       ��x���@�            �w@                           @1���~z@�            �u@������������������������       �>���2�@3            @U@������������������������       �V�� EE@�            0p@                           @r����@=           �@                          �9@C�[��_	@�           t�@                          �6@��~yC�@i           �@������������������������       ����}��@m            @e@������������������������       ��wv���@�            �y@                           �?�T��FA	@I           ؀@������������������������       ��:���@W            @a@������������������������       �[v�}m	@�            y@                           �?��6��d@�           0�@                           @���|@�            0r@������������������������       ���n@T             `@������������������������       ��9х?@h            `d@                          �:@�dm���@�            0t@������������������������       ���x�(s@�            �m@������������������������       ��a�as@;            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     ps@     �@      8@      J@     �{@     �U@     �@     �l@     ��@      w@      9@      @     �]@     �t@       @      2@      i@      <@     ��@     �V@     �~@     �c@      (@      @     �T@      h@      @      $@     �a@      0@     `o@     @R@     �j@     �W@      @              >@      J@              @      <@      �?     �^@      1@     �U@      <@      �?              $@      6@               @      .@      �?      N@      $@     �C@      $@      �?              4@      >@              �?      *@              O@      @      H@      2@              @     �J@     �a@      @      @      \@      .@      `@      L@     �_@     �P@      @      @     �G@     �V@      @      @     @T@      &@     �Q@      A@     �T@     �H@      @              @      I@       @       @      ?@      @     �M@      6@     �F@      1@                      B@     �`@      �?       @     �N@      (@     �}@      1@     `q@      P@      @              9@     @S@              @      B@       @     v@      (@     `h@     �C@       @              $@      9@              @      0@       @     �j@      @     �R@      0@       @              .@      J@               @      4@             `a@      @     @^@      7@                      &@      M@      �?       @      9@      $@     �]@      @     �T@      9@      @               @      8@                       @      @      5@      @      ,@      @      @              "@      A@      �?       @      1@      @     �X@             @Q@      5@       @      $@      h@     �j@      0@      A@     `n@     �M@     0s@     �a@     @r@     �j@      *@       @     `b@     @a@      &@      9@     �d@      H@     �b@     �]@      a@     �c@      (@      �?     @W@     �R@       @      .@      X@      ,@     @W@      G@     @R@      L@       @      �?     �B@      ;@              @      1@       @      9@      3@      6@      ,@                      L@      H@       @      "@     �S@      (@      Q@      ;@     �I@      E@       @      @      K@     �O@      @      $@     @Q@      A@     �L@      R@     �O@     �Y@      @              &@      2@              @      3@              6@      *@      6@      <@              @     �E@     �F@      @      @      I@      A@     �A@     �M@     �D@     �R@      @       @     �F@     �R@      @      "@     �S@      &@     �c@      6@     �c@     �J@      �?       @      8@      F@      @       @     �E@      �?      S@      @     �N@      6@      �?       @      .@      "@               @      3@              A@              @@      ,@      �?              "@     �A@      @      @      8@      �?      E@      @      =@       @                      5@      ?@      �?      �?     �A@      $@     @T@      1@     �W@      ?@                      &@      6@      �?              2@       @     @R@       @     �Q@      9@                      $@      "@              �?      1@       @       @      "@      8@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@�{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �5@G١:xB@�	           ��@       	                    @�ެ\z@e           ��@                           �?�(c�@�           ��@                          �2@���$q@�            �w@������������������������       ��� �Cd@y            `g@������������������������       ��Ȥ��@v             h@                           �?�U�C�@�           (�@������������������������       �Υ����@�            @p@������������������������       �@>;��@6           ~@
                          �4@_x9Q�@�           d�@                           �?$����l@@           X�@������������������������       ��tW��/�?�            �u@������������������������       ���I��@b           ��@                            �?��	���@`            �a@������������������������       ���|�^@3            �R@������������������������       ��O���?-            �P@                           @����A�@E           <�@                           �?����o	@�           ��@                           �?4��=@�            �q@������������������������       �V;;�o@P             ^@������������������������       �2����@q            @d@                           �?�2Fc��	@            (�@������������������������       �U1���?@�            0r@������������������������       ��I:��	@V           �@                           @r��@�           ��@                           �?8�$>�@{           ��@������������������������       �2(���'@p            �e@������������������������       ��M�T7@           y@������������������������       ���Ԭ�?	             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@     ps@     8�@      >@      O@     {@      R@     �@     �k@     ��@     �v@      :@      "@     �]@     `s@      .@      5@     @i@      8@     ��@     @T@      ~@     �e@      &@      "@      U@      e@      &@      ,@     �b@      2@     �p@     �P@     �i@     @^@      "@              =@     �I@       @      @      C@      @      `@      (@     @U@      ;@      �?               @      ;@                      :@       @     @P@      @     �F@      &@                      5@      8@       @      @      (@      �?     �O@      "@      D@      0@      �?      "@     �K@     @]@      "@      $@     @\@      .@      a@      K@     @^@     �W@       @      @      8@      I@       @      @      C@      "@      E@      3@      6@      D@      �?      @      ?@     �P@      �?      @     �R@      @     �W@     �A@     �X@      K@      @             �A@     �a@      @      @     �I@      @     �|@      .@     @q@     �I@       @             �@@     @^@      @      @     �D@      �?     z@      ,@      l@     �G@                      *@     �A@              �?      (@             �h@      @      Q@      ,@                      4@     �U@      @      @      =@      �?     @k@      $@     �c@     �@@                       @      5@               @      $@      @     �E@      �?      J@      @       @              �?      1@               @      @      @      .@      �?      ;@      �?                      �?      @                      @              <@              9@      @       @      &@      h@      n@      .@     �D@     �l@      H@      s@     �a@     �s@     �g@      .@      $@      b@     �d@      &@     �A@     �d@     �B@     �`@     @\@     �e@     @b@      .@       @      8@     �G@       @      @     �H@      @      I@      *@     �F@     �B@      @      �?      "@      3@               @     �@@      @      2@      @      0@      (@      @      �?      .@      <@       @      @      0@       @      @@      "@      =@      9@               @     @^@     �]@      "@      >@     @]@      @@     @U@      Y@     �_@     @[@      (@              >@      G@              3@     �B@      @      C@      4@      O@      ?@      @       @     �V@     @R@      "@      &@      T@      =@     �G@      T@     @P@     �S@      @      �?     �G@     �R@      @      @     @P@      &@     `e@      <@     �a@      E@              �?     �D@     �R@      @      @     �M@      &@     `e@      8@     �a@      E@                      @      >@                      *@      @      P@      @      F@      @              �?     �B@     �F@      @      @      G@      @     �Z@      1@     �X@     �B@                      @              �?              @                      @                        �t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJճ�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @%Y��@@�	           ��@       	                   �2@A��rl�@z           T�@                           @�=x��@A           H�@                           �?�+��G@�            �y@������������������������       �_)�@]            `b@������������������������       �߆�J[�@�            �p@                          �0@��}�@F            �[@������������������������       ��c�@�� @             =@������������������������       �벮<
�@8            @T@
                           �?iд)5U	@9           ��@                            @iX��@�           @�@������������������������       �m@+	�>@           0z@������������������������       ���R`	@�            �l@                          �4@A�m��d	@�           d�@������������������������       ��q-z@�            @m@������������������������       �x�Ȇf	@�           x�@                           @{s<�V�@(           |�@                           �?*j�Y	@�           �@                           @�f	BT��?�             v@������������������������       �2�a���@R            �_@������������������������       �������?�            �l@                          �7@F�)$L@�           Ȉ@������������������������       �m��@�           8�@������������������������       �}�K�p�@u            @f@                          �>@�P,@I            �@                            �?q���^�@<           x�@������������������������       �|�X��@K             `@������������������������       ��Q�/@�            �x@������������������������       �B�����@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        6@     �r@     0�@      D@      D@     �|@     @R@     ��@     `k@     p�@     Pu@     �A@      4@     �l@     �s@      <@      >@     �s@      N@     �x@     @g@     �w@     �l@      ;@      @      E@     �P@              @     �Q@      �?     �c@      B@     �X@     �D@       @       @     �@@     �G@               @      I@      �?     �_@      ;@     �V@      ?@               @      *@      3@                      ;@      �?      E@      &@      9@      @                      4@      <@               @      7@             @U@      0@     �P@      8@               @      "@      4@              �?      4@              =@      "@       @      $@       @               @      $@                       @              &@       @               @               @      @      $@              �?      2@              2@      @       @       @       @      0@     �g@      o@      <@      ;@     `n@     �M@      n@     �b@     �q@     �g@      9@      @      K@      ]@      &@      @     �V@      9@      Y@     �Q@     �V@     @R@      "@              ;@     @R@      @       @     �J@      .@      S@      M@      M@      G@      @      @      ;@     �E@      @      @      C@      $@      8@      (@      @@      ;@      @      *@     �`@     �`@      1@      5@      c@      A@     �a@      T@     �g@     @]@      0@      @      4@      2@      @      @      B@      @     �B@      &@      O@      :@      @      "@     �\@     �\@      &@      2@      ]@      >@      Z@     @Q@      `@     �V@      "@       @      R@     @m@      (@      $@     �a@      *@     x�@     �@@     0{@     �[@       @       @     �D@     �c@      @      @     �V@       @     �|@      1@      r@      Q@      @              $@      G@                      (@      @      h@      @     @S@      "@                      @      6@                      @       @     �I@       @     �@@      @                      @      8@                       @      �?     �a@       @      F@      @               @      ?@     @\@      @      @     �S@      @     �p@      *@     `j@     �M@      @              2@     �Y@      @       @      L@      @     `k@      &@     �c@      A@      @       @      *@      &@              �?      6@              G@       @     �J@      9@      @              ?@     �R@      @      @     �J@      @     �d@      0@     `b@      E@      �?              ;@     �R@      @      @     �I@      @     �d@      .@      b@      A@      �?              @      @      �?      �?      &@      �?      M@      @      A@      @                      7@     �P@      @      @      D@       @     �Z@      &@     �[@      ;@      �?              @      �?      �?               @       @              �?       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���ZhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��]�l@�	           ��@       	                    �?{�w-\�@           ƥ@                           �?�t�{	@X           ��@                          �<@�a��,	@�            `t@������������������������       �R�}[4�@�            �q@������������������������       �r��?
@            �D@                           �?s��aY	@�           X�@������������������������       �)���|@f            �d@������������������������       �wvT�
@"           `z@
                           @6S)��@�           H�@                          �1@�gZ���@�           ��@������������������������       ���c�|��?�             x@������������������������       ��sř��@�           ��@                           @���4(�@             D@������������������������       �ܢ]�1�@             =@������������������������       ��� 8��@             &@                           @�RD�=O@�           ��@                          �3@���9�	@           Ȋ@                          �2@�V���d@�            q@������������������������       �e����@z             i@������������������������       ���A=�@-             R@                          �:@�����%	@h           @�@������������������������       ���2v�@           @z@������������������������       �\iG��1
@f            �d@                          �9@u��@�            �p@                           @�m�b9@�            �k@������������������������       �߭�8�m @D            @\@������������������������       ���E@H            �Z@                           @]*#�`l@            �H@������������������������       �`��3I�@             9@������������������������       ��[����?             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      r@     ��@      B@     �G@     p{@     �X@     @�@     `n@      �@     �u@      =@      "@     �i@     �x@      2@      8@     �r@     �Q@     X�@     �e@     x�@     �l@      5@      "@      Y@      a@      &@      (@     @\@     �E@     @^@     @X@      b@     @[@      0@       @      <@      N@      @       @      C@      6@     �F@      H@      B@     �A@      @       @      8@      L@      @       @      C@      ,@     �E@     �D@      A@      5@      @              @      @                               @       @      @       @      ,@              @      R@     @S@       @      $@     �R@      5@      S@     �H@     @[@     �R@      "@              2@      9@                      ;@              @@      @     �E@      (@      @      @      K@      J@       @      $@      H@      5@      F@      F@     �P@      O@      @             @Z@     Pp@      @      (@     @g@      ;@     ��@     �S@     �{@     @^@      @             @Y@     @p@      @      (@     �f@      5@     p�@     �P@     `{@      ^@      @              @     �A@              @      1@             �h@      &@     @Y@      2@                     �X@      l@      @      "@     �d@      5@     �z@     �K@     u@     �Y@      @              @      �?      �?              @      @      @      (@       @      �?                       @      �?      �?                      @      @      (@      @      �?                       @                              @       @      �?              @                      &@     @U@     @d@      2@      7@     �a@      <@     �o@      Q@     �j@     @]@       @      &@     �R@     �`@      (@      4@     �_@      9@     �c@     �O@     ``@      X@       @      @      *@     �C@              $@      4@      @     �S@      ,@      I@     �A@      @      @      "@      ?@              @      4@              N@      (@     �B@      7@              �?      @       @              @              @      2@       @      *@      (@      @      @     �N@     @W@      (@      $@     �Z@      3@     @T@     �H@     @T@     �N@      @      �?     �@@      S@      @      @     @U@      &@     @P@      >@     @Q@      A@      @      @      <@      1@      @      @      5@       @      0@      3@      (@      ;@       @              &@      >@      @      @      ,@      @     �W@      @     �T@      5@                      &@      >@      @       @      @      @      T@       @      P@      2@                      @      ,@                       @      �?     �E@      �?      E@      @                      @      0@      @       @      @       @     �B@      �?      6@      ,@                                      @      �?      @              ,@      @      2@      @                                              �?      @              @      @      @       @                                      @                               @              (@      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJV�KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @6�[@�	           ��@       	                    �?�:�j+�@~           ��@                          �8@'�,�=	@            �@                           @��.nb@�           ؑ@������������������������       ���i��@�           (�@������������������������       ��.Q�Z�	@           {@                           @����m
@B           ��@������������������������       �hP�(V�	@           @}@������������������������       �6�r
e�	@(             O@
                           �?/$4�Q-@v           ��@                          �<@ ;��@|             g@������������������������       ���'��@t            �e@������������������������       ���q`�@             &@                           �?�(4�@�            `x@������������������������       ��"X�G@d            �b@������������������������       �	�PNuK@�             n@                          �7@��U�@0           �@                           �?�Ee�|@9           ��@                            @������?4           `~@������������������������       ����䨗�?           �y@������������������������       �rI��
�?3            �S@                           @�%�=�@           Ȉ@������������������������       ��P�l*@~            �g@������������������������       ��`����@�           �@                           �?�=<�-@�            @x@                            �?jf#2�� @<            �U@������������������������       �gx��� @             7@������������������������       �caRg�;�?.            �O@                          �<@ �^�a�@�            �r@������������������������       �VD7���@�            �n@������������������������       �y�8�=@$             M@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �r@     Ё@      ;@      J@     0|@     @T@     ��@     �k@     �@     0u@      B@      6@      l@     �t@      4@      E@     �s@      N@     �u@      g@     0z@     @o@      ?@      6@     �f@     �p@      3@     �A@     `l@     �E@     �j@     �a@     pr@      i@      ;@      @     �\@      g@      *@      6@     �c@      2@     �f@     �S@     �l@     @^@      ,@      �?     �P@     �Z@      @      $@     �W@      @      b@      B@     �c@     �S@      @      @      H@     �S@      @      (@      P@      .@      C@      E@      R@     �E@      "@      .@     �P@     �T@      @      *@     @Q@      9@      ?@      P@     @P@      T@      *@      @      N@     �R@      @      *@     �N@      4@      <@     �I@     �N@     @S@      $@       @      @      @      �?               @      @      @      *@      @      @      @             �E@      Q@      �?      @     �U@      1@     �`@     �E@      _@     �H@      @              &@      0@              �?      5@      @     @P@       @     �I@      *@      �?              &@      .@              �?      0@      @      P@              I@      *@                              �?                      @              �?       @      �?              �?              @@      J@      �?      @     @P@      ,@     �P@     �D@     @R@      B@      @              @      2@      �?      @      7@      @      4@      3@      ?@      4@      @              9@      A@               @      E@      &@     �G@      6@      E@      0@               @     @S@     `m@      @      $@     @a@      5@     ��@     �B@     �y@     @V@      @              M@     �h@      @      @     �T@      1@     �@      0@     �r@     �G@      @              2@     �P@               @      :@             �p@      @      W@      $@                      0@     �O@              �?      7@             `k@      @      R@      $@                       @      @              �?      @             �H@              4@                              D@     �`@      @       @      L@      1@     Pq@      (@     @j@     �B@      @              2@      D@                      @      *@      O@      @      >@      &@      @              6@     @W@      @       @     �H@      @     �j@       @     �f@      :@      �?       @      3@      B@       @      @      L@      @     �U@      5@      \@      E@      �?                      ,@                      @              ?@      @      =@      @                                                       @               @      @       @      �?                              ,@                      �?              7@       @      5@       @               @      3@      6@       @      @     �J@      @      L@      .@     �T@     �C@      �?       @      .@      2@      �?      @     �A@      @     �J@      ,@     �P@      =@      �?              @      @      �?      �?      2@              @      �?      0@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$[�EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?3�~� M@�	           ��@       	                    @���3�@            L�@                          �9@�$a�f@�           ��@                           �?��G�Ԍ@K           P@������������������������       �2����@�            �m@������������������������       �� �,�@�            �p@                           �?����B�@\             `@������������������������       �x�"�@)             L@������������������������       ����\@3            @R@
                          �8@f��38@Y           �@                           @}���'� @*           p}@������������������������       ��D!��7�?�            ps@������������������������       ��#<�!�@i             d@                          �:@�Sw��@/            �Q@������������������������       �R(H��4�?             :@������������������������       �^��}��@             F@                           �?Y��׍@�           l�@                           �?��B��	@�           �@                           @�c��F@           P{@������������������������       ��q��w�@8            �T@������������������������       �,(��@�             v@                            @<>���	@�           8�@������������������������       �$S��	@�            pw@������������������������       ��LoY �	@�             u@                           @_�)��@�           �@                          �5@c�U�`@W           t�@������������������������       �K=_���@           ��@������������������������       ��<��:X@S           (�@                           !@滉*@|            �k@������������������������       ���/�j@q            �h@������������������������       �o�*��@             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      q@     ��@      7@      N@     �}@      S@     ��@     �k@     `�@      w@      B@      @      Q@     �d@       @       @     @X@      &@     �x@     �D@     0r@     �S@      @      @     �L@     �S@              @     �Q@      @      b@     �A@      e@     �L@      @             �G@      K@              @      F@      @      `@      7@     `b@     �E@      @              6@      3@              @      :@      @     @R@      (@     �J@      6@       @              9@     �A@               @      2@              L@      &@     �W@      5@       @      @      $@      8@              �?      :@      �?      0@      (@      5@      ,@      �?      @      @       @                      "@      �?       @       @      "@      @                      @      0@              �?      1@               @      @      (@      @      �?              &@     @V@       @      �?      ;@      @     �o@      @     �^@      6@      �?              &@     �S@       @      �?      9@      @      m@       @      Y@      .@      �?              @     �G@                      *@      @      e@      �?      P@      @                      @      ?@       @      �?      (@              P@      �?      B@       @      �?                      &@                       @      @      4@      @      7@      @                              �?                              @      @              *@      @                              $@                       @              ,@      @      $@      @              .@     �i@     �x@      5@      J@     �w@     @P@     P�@     �f@     H�@     0r@      >@      (@     @]@     �d@      ,@      @@      j@      E@     @_@     �Z@     �c@     �b@      5@      �?      A@     �N@       @      .@     �T@      $@     �R@      =@     @R@     �I@      @      �?      @      &@               @      1@      @      @      @      4@      @                      ;@      I@       @      *@     @P@      @     @Q@      7@     �J@      F@      @      &@     �T@     �Y@      (@      1@     �_@      @@      I@     �S@     �T@     �X@      1@      @      I@     �E@      @      "@      O@      1@      ;@     �J@     �A@      N@      @      @     �@@      N@      @       @     @P@      .@      7@      9@      H@      C@      $@      @     �U@     `m@      @      4@     �d@      7@     �|@     �R@     �v@     �a@      "@      @     @P@     �i@      @      3@     �b@      3@     Py@      J@     @u@      \@                      6@      b@      �?      $@      R@      @     �r@      7@     �k@      M@              @     �E@      O@      @      "@      S@      (@     @[@      =@     @]@      K@                      6@      =@      @      �?      3@      @      L@      7@      9@      >@      "@              *@      :@      @      �?      ,@      �?      L@      6@      9@      =@      "@              "@      @                      @      @              �?              �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�(1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��8>�+@�	           ��@       	                     @�:�xU�@�           ��@                          �:@����0�@w           <�@                          �4@�طip@�           �@������������������������       �k�_�+C@\           �@������������������������       �n���	@}           ��@                          �=@W�ke@�            `q@������������������������       ����0y@^             e@������������������������       �|��W�@@            �[@
                           �?���$�?@           `�@                           �?,0>��@�           p�@������������������������       �V��/@|            �g@������������������������       �:��c��@4            @                          �3@��䒑�@k            �c@������������������������       �quQ�4 @'            �J@������������������������       �)���e@D            @Z@                          �1@�nd�J�@           ��@                            �?�n�V&�?�            �u@                           @m{7�?.            �S@������������������������       �4[�ji��?             I@������������������������       ���ē�q�?             =@                          �0@�����?�             q@������������������������       �}!4�]��?;            @Y@������������������������       �2c�S�g�?o            `e@                           @&ɉW�@A           <�@                           @<��	��@=           ��@������������������������       ������@j           ��@������������������������       ��&b�� @�            @u@                           �?X!�cI1@           �y@������������������������       �1�s�;�@�            �j@������������������������       �ͮ��=@            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     ps@     ��@      :@     �D@     �~@     �S@     Ȏ@     �j@     ��@     �v@      :@      .@     `l@     �u@      0@     �A@     Pv@      O@     @w@     `f@     �w@      p@      8@      $@      b@      h@      "@      3@     `l@      E@     �k@     �`@     �n@     �c@      1@       @     �^@      e@      @      2@     �d@      >@     �h@     �W@     �j@     �[@      *@      @     �C@      V@      @      @     �T@      @     �[@     �H@     �Z@      J@       @      @      U@      T@       @      .@     @T@      8@      V@      G@     �Z@      M@      &@       @      6@      9@      @      �?     �O@      (@      8@      C@      A@     �H@      @       @       @      4@      @      �?     �D@      @      ,@      0@      7@     �A@                      ,@      @                      6@       @      $@      6@      &@      ,@      @      @     �T@     `c@      @      0@     @`@      4@     �b@      G@      `@     @X@      @      @     @R@     �_@      @      ,@     �\@      1@     �X@     �D@     �Z@     �S@      @              2@      B@              @      :@      @     �I@      @      >@      *@              @     �K@     �V@      @      $@     @V@      ,@     �G@      A@      S@     @P@      @              "@      =@      �?       @      .@      @      J@      @      7@      3@                      �?      @               @                      <@      @      $@       @                       @      6@      �?              .@      @      8@       @      *@      1@                      U@      l@      $@      @     �`@      1@     (�@     �A@     �y@     �[@       @              @     �B@              �?      ,@             �g@       @      U@      .@      �?                      @              �?       @              J@      �?      (@      @                              @                      �?             �A@              @      @                               @              �?      �?              1@      �?      @                              @      @@                      (@             `a@      �?      R@      "@      �?                      4@                       @              L@              4@      @                      @      (@                      $@             �T@      �?      J@      @      �?             �S@     `g@      $@      @     �]@      1@     `z@     �@@     �t@     �W@      �?             �E@      a@       @      @     �S@      $@     Ps@      1@     �l@      J@      �?             �B@      R@       @             �K@      $@     �e@      .@      a@      E@      �?              @     @P@              @      7@              a@       @     �W@      $@                     �A@      I@       @       @     �D@      @     @\@      0@     �X@     �E@                      1@      :@      @       @      8@      @      P@      @      G@      6@                      2@      8@      @              1@      @     �H@      "@      J@      5@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ
Դ1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�w"�GX@�	           ��@       	                   �2@���Zc�@�           ~�@                           �?����p�@2           �@                          �1@�uE�]�@z            �j@������������������������       �=�!YI�@E            �]@������������������������       ��M:b�a@5            @W@                           @�ARS*�@�            �r@������������������������       �	��)��@�             n@������������������������       � W�>�@!             L@
                           �?^� N	@b           �@                           �?)f�q�@1           �}@������������������������       �>�����@�            �v@������������������������       ����]J@M             \@                           @�=���	@1           ��@������������������������       �"X%��	@�           ̐@������������������������       �!�$8@n            �f@                          �4@��F�@6           (�@                           �?=��H�s@E           @�@                          �1@�h��K;�?�            0u@������������������������       �N�(h� �?_             c@������������������������       �����FL�?y            @g@                           �?n�&N_C@m           ��@������������������������       �	kV�]@�            0r@������������������������       �6("s�@�             q@                          �7@x���)@�           �@                           @ᖃ�0@�            `w@������������������������       �`��7�@�            `p@������������������������       �r j�s"@J             \@                          �<@�=��D|@           �x@������������������������       ���nT@�            �r@������������������������       ��4��/�@;            �W@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     �@      :@     �N@     �{@     �V@     (�@     �m@     �@     pw@      ;@      0@     �i@     Pt@      4@     �D@     �t@     @R@     pw@     `h@      x@     p@      5@      �?      ;@     �T@              @     �P@      @     @a@     �B@     @[@     �A@              �?      "@     �@@                      >@      @     �P@      7@      @@      .@                      @      3@                      &@      �?      D@      4@      .@      $@              �?      @      ,@                      3@       @      :@      @      1@      @                      2@      I@              @     �B@      @      R@      ,@     @S@      4@                      ,@      @@              @      <@              N@      &@     �Q@      4@                      @      2@              �?      "@      @      (@      @      @                      .@      f@     @n@      4@      B@     Pp@     �P@     �m@     �c@     0q@     �k@      5@      �?      M@     �J@              @     �J@      @     @[@     �@@      Z@     �I@      @      �?      H@     �D@              @     �G@       @     @R@      <@     �R@     �E@       @              $@      (@                      @       @      B@      @      =@       @      @      ,@     �]@     �g@      4@     �@@      j@     �O@      `@     @_@     `e@     `e@      .@       @     @X@     `d@      4@      @@     �e@     �L@      \@      V@     �d@     �b@      (@      @      6@      :@              �?      A@      @      0@     �B@      @      7@      @      �?     @T@     �k@      @      4@     �\@      2@     ��@      F@      x@     �]@      @             �@@     �X@      @      $@     �C@      @     �{@      0@     �j@      G@      �?              "@      >@              @      .@              h@      @     �Q@      $@      �?              @      $@              @      $@             �V@              ;@      @      �?              @      4@              �?      @             �Y@      @      F@      @                      8@      Q@      @      @      8@      @      o@      &@     �a@      B@                       @      8@      @       @      3@      �?     �_@       @     @S@      6@                      0@      F@               @      @      @     @^@      @     �P@      ,@              �?      H@     �^@      @      $@      S@      ,@     `k@      <@     �e@      R@      @              3@      R@      @      @     �@@      "@     �_@      @     @R@      :@      @              2@      H@                      5@      @     @Y@      @     �G@      .@      @              �?      8@      @      @      (@      @      9@       @      :@      &@              �?      =@      I@              @     �E@      @     @W@      7@     �X@      G@       @      �?      2@      ?@              @      9@      @      S@      0@     �U@     �B@       @              &@      3@                      2@              1@      @      *@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��8!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�pam@�	           ��@       	                    �?�6
@           ��@                          �7@�=�'>@A           ��@                           �?k�����@�           ��@������������������������       �a�ZNq@�             w@������������������������       ��l���e@�             t@                           �?�Uo@�@�            `l@������������������������       ����i[@>            �Y@������������������������       ���yW2�@Q            @_@
                           �?�OW)�@�           ��@                           �?��~�@�            �@������������������������       ���&���@�            �h@������������������������       ��S����@h           �@                           �?t���o�@�           ��@������������������������       ��)M�ۯ	@8            �X@������������������������       ���C��}@�           �@                           �?����I@�           (�@                           �? BHi-@�            �r@                          �7@N�?Wn�@m            �e@������������������������       �.`R��@I             ^@������������������������       �uG�(M�@$             J@                           �?41�L4��?[             `@������������������������       �b��o� @/            �Q@������������������������       ���e��?,            �M@                           �?B��@�@�           �@                           �?g��Z��	@@           �@������������������������       �f�`4��@`             b@������������������������       �8�	@�            �v@                           @|����@�            @r@������������������������       �H����@�            `p@������������������������       �����X@             >@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ?@     �r@     ��@      B@      G@     `z@     �U@     ��@     `j@     �@     �v@      A@      (@     �i@      y@      2@     �D@     r@     @P@     ��@     �b@     ��@     @o@      7@       @     �K@      a@              @     @P@      *@     �s@      2@     `m@      M@      @              A@     @Y@              @      K@      @     �q@      $@     �d@      @@      �?              *@      J@              @     �B@      @     �d@      @     �R@      $@                      5@     �H@                      1@             �\@      @      W@      6@      �?       @      5@      B@              �?      &@       @     �C@       @     @Q@      :@      @       @      .@      4@              �?      @       @      @      @      ;@      ,@      @              @      0@                      @      @      @@      @      E@      (@       @      $@     �b@     �p@      2@     �A@      l@      J@     �y@     ``@     �x@      h@      0@             @P@     �\@       @      1@     �W@      .@     �e@      I@     @b@     �R@      ,@              1@     �E@      @       @      6@       @      ;@      <@      (@      ;@      $@              H@      R@      @      .@     @R@      @      b@      6@     �`@      H@      @      $@     �U@     �b@      $@      2@      `@     �B@      n@     @T@     �n@     @]@       @      @      @      &@              "@      *@      @      0@      $@      0@      @              @     @T@     `a@      $@      "@      ]@      >@      l@     �Q@     �l@     �[@       @      3@     @W@     �d@      2@      @     �`@      6@     0p@      O@      i@     �[@      &@              :@     �B@       @      �?      @@             �Y@      "@      R@      3@                      4@      A@       @      �?      6@              C@      @      A@      ,@                      &@      9@                      @              ?@      @      @@      (@                      "@      "@       @      �?      0@              @      @       @       @                      @      @                      $@             @P@       @      C@      @                      @      �?                       @             �@@              2@      @                      �?       @                       @              @@       @      4@                      3@     �P@     �_@      0@      @     @Y@      6@     �c@     �J@      `@      W@      &@      3@      J@      T@      (@      @     @R@      4@      O@      E@     @R@      N@      "@      @      .@      6@      @       @      5@      �?      <@      $@      4@      0@      @      0@     �B@      M@      "@      �?      J@      3@      A@      @@     �J@      F@      @              .@     �G@      @      �?      <@       @     �W@      &@      L@      @@       @              $@      C@      @      �?      6@       @     �V@      $@     �J@      @@                      @      "@      �?              @              @      �?      @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ�~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�<�J�@�	           ��@       	                   �1@5튞�.@�           ��@                          �0@��٪iQ�?�            �p@                           �?~�Vb/��?7            �V@������������������������       ��+P&� @            �F@������������������������       ��[��$�?             G@                           @�M����?i            @f@������������������������       �"S�����?Q            @a@������������������������       ��1��\�?             D@
                           �?Y����-@H           ��@                          �8@������@�            �v@������������������������       ��x(���@�            @o@������������������������       �GLd-@O            �\@                            @��5pj�@b           ��@������������������������       ���> .7@&           �}@������������������������       ��q�٨G�?<            @U@                           @T�ދ�@�           :�@                           �?�ቦ��	@�           T�@                          �:@�4�[�

@�           ��@������������������������       �X�!�Ŭ	@6           Ћ@������������������������       ��N�;�	@�            �n@                          �5@�m�{e@           `z@������������������������       ����~@�            �l@������������������������       �P'�ƨZ@u             h@                          �7@���@�            �@                           �?erc�+@           Љ@������������������������       ��%��D@#             K@������������������������       �Q�d��@�            �@                           @��h2@�            �t@������������������������       ��!�	;z@�            p@������������������������       ��s�5L@)            @S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     Ps@     h�@      ?@     �Q@     P|@     �W@     0�@     �i@     ��@     �v@      B@             �S@     �d@       @      $@     @V@      1@      }@      >@     `p@     �Q@       @              @      ;@                      8@             `d@      @      C@      @                      �?      (@                      0@              H@      �?      "@      @                              @                      $@              5@      �?      @      �?                      �?      @                      @              ;@               @      @                      @      .@                       @             �\@      @      =@       @                       @      ,@                       @             �W@      @      4@       @                       @      �?                      @              4@       @      "@                             @R@     `a@       @      $@     @P@      1@     �r@      8@      l@      P@       @              H@      N@              @     �B@      �?     @P@      2@     @V@     �@@       @             �@@     �A@               @      0@      �?      M@      $@      R@      1@      @              .@      9@              @      5@              @       @      1@      0@       @              9@     �S@       @      @      <@      0@     �m@      @     �`@      ?@                      5@     �R@       @       @      9@      0@     �g@      @     �\@      <@                      @      @               @      @             �G@      �?      4@      @              9@     �l@     pv@      =@     �N@     �v@     @S@     ��@      f@      @     �r@      <@      9@     �c@     @k@      4@     �F@     `o@     �M@     `i@     �a@     �k@     �g@      :@      9@     �^@      c@      3@      =@     �h@      G@     `a@     �V@     �a@     `b@      8@      ,@     �X@     �`@      "@      8@     �c@      B@     �\@     @P@      `@     �V@      4@      &@      9@      5@      $@      @     �C@      $@      9@      9@      ,@      L@      @              B@     @P@      �?      0@      K@      *@      P@     �I@     �S@     �D@       @               @      D@      �?      &@      <@      @      H@      8@     �D@      8@                      <@      9@              @      :@       @      0@      ;@      C@      1@       @              R@     �a@      "@      0@     @\@      2@     w@      B@     @q@      [@       @             �B@     @Z@       @       @      M@      (@     �s@      1@     �h@     �P@       @              @      "@                       @      @      @      @      &@      @                      ?@      X@       @       @      I@      @     0s@      ,@     `g@      O@       @             �A@      B@      �?       @     �K@      @     �K@      3@     �S@     �D@                      0@      ;@               @      E@      @     �G@      (@      Q@     �@@                      3@      "@      �?              *@       @       @      @      $@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�|hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��o@�	           ��@       	                    �?&�sP�h	@           ��@                           �?/�H
 @/           �}@                            @|8��sM@t            �g@������������������������       ��蔎@U            �_@������������������������       ��f�V���?             O@                            @4}殹�@�            �q@������������������������       �yKԠ.@_            �a@������������������������       �Y�GĻ@\             b@
                            �?U,6 d�	@�           ��@                           @~��E9�@�            �v@������������������������       ��i�^�-@�            �j@������������������������       ���dޗ�@X            �b@                           @�d��b
@�           ��@������������������������       ��>u�(�	@�            �@������������������������       �H��/X�@             6@                           �?��O_p#@�           �@                            �?�`�&4�@�           �@                           @s�T�	 @u            �g@������������������������       ��/���f�?!             N@������������������������       ��O((�6�?T             `@                           @�}A9�=@c           0�@������������������������       �J[��o�@�            �k@������������������������       �l����� @�            pt@                           @@���F8@�           ��@                           �?���]@�           ��@������������������������       ��":�@            �F@������������������������       �����b@�           x�@                           �?���@+           X�@������������������������       ����C�@#             K@������������������������       �G����@           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     h�@      @@      L@     P{@     @R@     ��@      n@     Ї@     �v@     �A@      3@     @f@     `m@      7@      <@     �l@      G@     `m@     �b@     @m@      h@      ;@      �?     �K@     @S@      �?       @     �L@      @     �[@      >@     �V@      C@      @      �?      .@      :@                      5@             @P@      @      F@      "@      @      �?      *@      0@                      1@              =@      @      B@       @      @               @      $@                      @              B@      �?       @      �?                      D@     �I@      �?       @      B@      @      G@      9@      G@      =@       @              .@      0@      �?      @      5@       @      8@      "@      ;@      5@       @              9@     �A@              @      .@      �?      6@      0@      3@       @              2@     �^@     �c@      6@      4@     �e@     �E@      _@      ^@      b@     `c@      6@      @      G@     �C@       @      @      P@      @     �H@     �L@     �B@     �G@      $@      @      7@      <@      �?              D@      @      9@      =@      8@      A@       @              7@      &@      �?      @      8@      �?      8@      <@      *@      *@       @      .@     @S@     �]@      4@      .@     �[@     �B@     �R@     �O@     �Z@      [@      (@      (@     @S@     @]@      4@      .@     @Z@      B@     �R@     �M@     �Z@     @Z@      "@      @               @                      @      �?      �?      @              @      @       @     @a@      t@      "@      <@     �i@      ;@     ��@     �V@     ��@     �d@       @              8@     �X@       @      @     �B@      &@     �u@      *@     `e@     �@@      �?              �?      ;@       @       @      "@      @     @X@             �E@      @                      �?      @               @              �?      :@              7@                                      4@       @              "@      @     �Q@              4@      @                      7@      R@               @      <@      @     �n@      *@      `@      =@      �?              .@      >@                      .@      @      W@      @      E@      0@                       @      E@               @      *@             `c@      @     �U@      *@      �?       @     �\@     �k@      @      8@      e@      0@     �{@     �S@     Pv@     �`@      @       @     �Q@     �Z@              "@     �U@      &@     �c@     �J@     ``@      Q@      @       @       @      @               @      $@               @       @       @      $@                      O@      Y@              @      S@      &@     `c@     �I@      `@      M@      @              F@      ]@      @      .@     �T@      @     �q@      9@     @l@     �P@      �?                      @              �?       @              &@       @      6@      @                      F@      \@      @      ,@     @T@      @     @q@      1@     �i@      N@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJz��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��řj@�	           ��@       	                    �?MZ>N_	@           8�@                           �?+��(d@�           �@                          �1@�:�$@x            @h@������������������������       �N�+���?            �H@������������������������       �4NT���@]             b@                          �=@�T��L�@           �{@������������������������       �*�H�@           �y@������������������������       ��=f���@             @@
                            �?�$a��	@t           ��@                           �?M����@�            �r@������������������������       �)(����@3             W@������������������������       ���;X�@�             j@                           @�vNXy
@�           (�@������������������������       ��<�CV�	@�           @�@������������������������       ��]#l��@*            �N@                          �7@�ܱ�V@�           ��@                           �?-�A�y@9           ��@                           @%	�F� @v            �@������������������������       �Va/�C@�             q@������������������������       ��? ^F�?�             u@                           @+jϦ�G@�           �@������������������������       ���`S�5@*            @������������������������       ��flI�@�           ��@                            @���2@`           ��@                            �?2بET@            z@������������������������       ��z�I<�@�            �p@������������������������       �@y��@]            �b@                           @?"dڬ@R            @]@������������������������       �|���*n@;            �T@������������������������       ��� s�W@             A@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     x�@      =@     �N@     �}@     �T@     ��@     `i@     (�@     �v@      B@      4@     �f@     �n@      2@     �C@      n@      F@     �l@     @_@     @n@      i@      <@      �?     �K@     @Y@       @      .@     �W@      1@     �\@     �C@     �[@     �R@      *@      �?      4@      6@                      9@             �K@      @      H@      .@      @               @      �?                      (@              5@              &@       @              �?      2@      5@                      *@              A@      @     �B@      *@      @             �A@     �S@       @      .@     �Q@      1@      N@      A@      O@     �M@      $@              >@     �S@      �?      .@     �Q@      0@      L@      >@     �M@      G@      $@              @      �?      �?                      �?      @      @      @      *@              3@     �_@      b@      0@      8@      b@      ;@      ]@     �U@     �`@     �_@      .@             �G@      C@      �?      @     �C@       @     �C@      >@      D@      H@      @              0@      $@                      "@      �?      9@       @      *@      $@                      ?@      <@      �?      @      >@      @      ,@      6@      ;@      C@      @      3@      T@     �Z@      .@      1@     �Z@      3@     @S@      L@      W@     �S@      (@      .@     �S@     �X@      .@      1@     @W@      0@     @Q@      H@     �V@     @Q@      @      @       @      @                      *@      @       @       @       @      "@      @       @     @]@     �s@      &@      6@     @m@      C@     h�@     �S@     ��@     `d@       @             �Q@      p@      &@      .@     `e@      =@     �@      D@     �x@     @X@      @              2@     �S@       @      @     �G@      @     `s@      @     �_@      1@      �?              .@      B@              �?      <@      @     �]@      �?     �N@      "@                      @      E@       @       @      3@              h@      @     �P@       @      �?              J@     �f@      "@      (@      _@      8@     �v@      B@      q@      T@       @              8@     @W@      @      @     �L@      6@      b@      :@     �V@      >@      �?              <@     �U@      @       @     �P@       @     @k@      $@     �f@      I@      �?       @     �G@      L@              @     �O@      "@      [@      C@     �`@     �P@      @       @      >@      H@              @      H@      "@      S@      =@     �[@     �J@      @              8@      ?@              @      5@      @      H@      4@     @S@      B@      @       @      @      1@               @      ;@      @      <@      "@     �@@      1@       @              1@       @              �?      .@              @@      "@      6@      *@                      *@      @                      $@              <@      @      .@      @                      @       @              �?      @              @      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��AhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@=��`�@�	           ��@       	                    �?v�	![@q           Ȝ@                           @ǰ��@�           �@                          �1@Z���G�@�            �r@������������������������       ��8�@9            @W@������������������������       ���_�y@}            �i@                           �?�0�7�?�            �u@������������������������       �WȩK�?�            �k@������������������������       �����N��?X             _@
                           @_�[[@�           Ē@                           @����]!@i           ��@������������������������       �m�/�@A           ��@������������������������       ����gN�@(            �Q@                          �1@qp"$�G@t           ؂@������������������������       �(�v~`��?}            �i@������������������������       ���[�|@�            �x@                           �?QF�7��@)           .�@                          �<@	{)S�i@{            �@                          �;@�u� ��@C           P~@������������������������       ��p+�@2           �|@������������������������       �MɉՀ@             8@                           �?���25@8            �V@������������������������       ��!� 0@%            �M@������������������������       �(<�*��@             @@                           @�]g{Z	@�           \�@                          �<@~ff�f-	@&            �@������������������������       �� Q���@�           ��@������������������������       ��]~y�@�            �j@                            �?�?�<�@�            �j@������������������������       ��ͧ,y\@*            �P@������������������������       �D�b�Y�@^            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �s@     p�@      5@     �P@     {@     �Y@     h�@      m@      �@     `v@      :@      @      X@     `p@      &@      2@     �c@      6@     ��@     @U@      y@     �b@      @             �@@     �R@              @     �G@      @     �q@      5@     �a@      ;@       @              7@     �B@              @     �@@      @     �T@      2@     �R@      4@      �?              @       @                      1@              ?@       @      7@      �?                      2@      =@              @      0@      @     �I@      $@     �I@      3@      �?              $@     �B@              �?      ,@             `i@      @      Q@      @      �?              @      5@              �?      *@             �`@              D@      @                      @      0@                      �?             �Q@      @      <@       @      �?      @     �O@     �g@      &@      (@     @[@      2@     �u@      P@      p@     �^@      @      @     �C@     @X@      @      @     �T@      (@     �_@     �K@     �V@      R@      @      @      A@     �V@      @      @     �P@      @     �]@     �D@     �U@      O@       @      �?      @      @                      .@      @       @      ,@      @      $@      �?              8@     �V@      @      @      ;@      @     `k@      "@     �d@      I@                      �?      ?@               @      @             �V@      @     �N@      $@                      7@      N@      @      @      6@      @      `@      @     �Z@      D@              0@     `k@     �r@      $@      H@     Pq@     @T@     `w@     �b@     @w@      j@      5@      �?     �J@      T@               @     �P@      @     `c@      ;@      _@      I@      @      �?      G@     �Q@              @     �K@      @     @a@      4@      \@      <@       @              D@      Q@              @      K@      @     �`@      4@     �Z@      <@       @      �?      @      @                      �?      @      @              @                              @      "@              @      (@              1@      @      (@      6@       @              @      @              @      @              @      @      @      3@                      �?       @                      @              *@      �?      @      @       @      .@     �d@      k@      $@      D@     @j@     �R@     `k@     @^@      o@     �c@      1@       @     �a@     �f@      "@      C@     @e@     �N@     �f@     �W@     �m@      b@      ,@      @     @\@      c@      @      =@      b@     �I@      d@     �P@     @k@     �Y@      ,@      �?      =@      =@       @      "@      9@      $@      3@      ;@      3@      E@              @      8@      A@      �?       @      D@      *@     �C@      ;@      &@      ,@      @              "@      &@      �?              @       @       @      *@      @       @       @      @      .@      7@               @     �A@      &@      ?@      ,@      @      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJj�"!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @o��-)@�	           ��@       	                    �?��ҽq�@j           $�@                          �4@�z�7(	@�           ̘@                          �2@w�p�@~            �@������������������������       �h�����@�            pt@������������������������       ��~�S�@�            �q@                           �?��VG��	@s           ��@������������������������       ��@7x�@�            u@������������������������       �A
s�|
@�           �@
                           �?�r2@y           ��@                          �<@�g��u@o            �g@������������������������       ���i� �@h             f@������������������������       ���q`�@             &@                            �?B��|�@
           0z@������������������������       �p����@O             ^@������������������������       �9��o@�            �r@                           @�9 ���@I           ܚ@                          �1@����@�           В@                           �?�L�?�            �p@������������������������       ��� [	��?b            @d@������������������������       ��yh�J�?H            �Z@                           @A��@E           8�@������������������������       ���r=�6@�            �@������������������������       �L�P�,�@�            0r@                           �?�S�X�@Z           �@                           �?;Fʵ�;@�            �g@������������������������       �'��ߒ@M            �[@������������������������       �*��s̥ @8            �S@                            �?g.p�&f@�            Pt@������������������������       ����@w            �f@������������������������       �/�&5@^            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �q@     (�@     �@@     �K@      {@     �R@     X�@      i@     p�@     �w@      :@      4@     �i@     �u@      :@      A@     Pr@     �M@     �y@     �d@     �u@     �o@      8@      4@      d@      o@      5@      :@      l@      G@     �p@     �_@     �l@     �h@      6@      @     �L@     @Q@      @      @     �T@      *@     @c@      C@     �Y@      R@      @      @     �A@     �B@      �?      @     �H@       @     �W@      4@      I@      <@       @       @      6@      @@      @      �?     �@@      &@     �M@      2@     �J@      F@      @      ,@     �Y@     `f@      1@      5@     �a@     �@@      \@     @V@      `@      _@      1@      �?      9@      L@      �?      @     �P@      $@      I@      >@     �I@     �B@       @      *@     �S@     �^@      0@      ,@     �R@      7@      O@     �M@     @S@     �U@      .@              F@     �Y@      @       @     @Q@      *@     @b@     �C@      ^@     �M@       @              1@      4@                      $@      @     @P@       @     �H@      *@      �?              .@      4@                      $@      @      P@      @      H@      (@                       @                                              �?      @      �?      �?      �?              ;@     �T@      @       @     �M@       @     @T@      ?@     �Q@      G@      �?              @      :@               @      .@      @     �@@      @      $@      .@      �?              5@      L@      @      @      F@      @      H@      8@     �N@      ?@               @     @S@     �l@      @      5@     `a@      .@     Ѓ@     �A@     �z@     @_@       @       @      M@     �c@      �?      @     �U@      $@     `~@      2@     �r@     �S@                      @      ?@                      $@             @d@       @     �K@      @                      @      5@                      @              X@       @      @@      �?                              $@                      @             �P@              7@      @               @      K@     @_@      �?      @     @S@      $@     @t@      0@     �n@     �R@               @      2@     �V@              @     �I@      "@     �m@       @      f@      F@                      B@      A@      �?              :@      �?     �U@       @      Q@      >@                      3@     �R@      @      ,@      J@      @     �b@      1@     ``@      G@       @              �?      @@               @      *@              T@       @      H@      (@                      �?      1@               @      $@             �J@      �?      6@      @                              .@                      @              ;@      �?      :@      @                      2@     �E@      @      (@     �C@      @      Q@      .@     �T@      A@       @              &@      9@              @      0@       @     �@@      "@     �L@      6@                      @      2@      @      @      7@      @     �A@      @      :@      (@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�
#ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?%�9�+x@�	           ��@       	                    @�ȻXZ�@�           ؒ@                            @#H����@�           `�@                          �;@�)8ތ@           �y@������������������������       �5
VM@�             w@������������������������       ��QS���@             E@                           �?#1έH�@�             n@������������������������       �2���2@J            @\@������������������������       �$���#@K            �_@
                            �?���@e           P�@                          �6@J���A�?O            @^@������������������������       �n�W.���?<            @W@������������������������       ��e��� @             <@                            @6�!:n@           {@������������������������       ��,�x�@�            0u@������������������������       ��1���??            �W@                           @p0G��T@�           &�@                           �?�5n�	@�           �@                            �?�4MB�@           �z@������������������������       �3*LR��@V            `a@������������������������       ���F��!@�            @r@                          �5@�v-��	@�           \�@������������������������       ��3��AN	@T           ��@������������������������       �� ���	@s           ��@                          �9@MZݗ{�@�           4�@                          �1@�X�3@\           ��@������������������������       ��5
o{�?�            �i@������������������������       ��o��c@�           @�@                            @v6���@u            �f@������������������������       �(rQ�g�@[             b@������������������������       �`L�-�@             C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     s@     Ȁ@     �B@     �N@     �z@      X@     ��@     `j@     ��@     0x@      @@      �?     @W@     �c@      @      "@     �W@      ,@     `z@     �H@     �q@      T@       @      �?     �S@      W@      �?       @      R@       @     `b@      B@      c@      K@       @      �?      N@     �I@      �?       @     �B@       @      U@      5@     @[@      B@       @              J@      H@      �?       @      A@      @      U@      3@     �W@      :@       @      �?       @      @                      @      �?               @      ,@      $@                      2@     �D@              @     �A@             �O@      .@      F@      2@                      @      *@              @      4@              :@      @      8@      (@                      &@      <@               @      .@             �B@       @      4@      @                      .@     �P@       @      �?      7@      @     0q@      *@     �_@      :@                               @       @              $@      �?     �Q@              1@      (@                               @                      @              N@              $@      &@                                       @              @      �?      &@              @      �?                      .@      M@              �?      *@      @     �i@      *@     �[@      ,@                      *@      L@              �?      $@      @     �b@      (@     @T@      (@                       @       @                      @             �K@      �?      =@       @              *@     �j@     �w@      A@      J@     �t@     �T@     ��@     @d@     ��@     0s@      >@      &@     `a@     �m@      8@     �F@     �k@     �P@     @h@     `a@      m@     �i@      ;@       @      .@     �Q@      �?      7@     @Q@      (@      P@      ?@     �R@     �O@      @              @      .@              (@      8@      @      9@      0@      >@      @      �?       @      "@     �K@      �?      &@     �F@       @     �C@      .@      F@     �L@      @      "@      _@     �d@      7@      6@     �b@      K@     @`@      [@     �c@      b@      4@      @     �C@      V@      @      &@     �P@      <@     @U@      K@     @X@      K@       @      @     @U@     �S@      0@      &@      U@      :@     �F@      K@      O@     �V@      (@       @     @R@     �a@      $@      @      \@      0@     `w@      7@     �r@      Y@      @       @      H@      `@      @      @     �T@      *@     �u@      *@     �o@     @T@      @               @      8@                      (@             �W@             �O@      @               @      D@     @Z@      @      @     �Q@      *@     �o@      *@     �g@     �R@      @              9@      *@      @       @      >@      @      :@      $@     �I@      3@                      8@      &@       @      �?      6@      @      0@      @     �D@      1@                      �?       @      �?      �?       @              $@      @      $@       @        �t�bub�N      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�s��*X@�	           ��@       	                    �?�)B�)@           T�@                          �8@�!	}��@3           0~@                           �?�;��(@�            �v@������������������������       �x�xw�@S            �_@������������������������       � ���+,@�            �m@                           �?��ؔ�@K            �]@������������������������       �Iٗ�j@             B@������������������������       ��(��@2            �T@
                           @;zf@�           ��@                          �3@;�%m@t            �g@������������������������       �Nj��U@2            �R@������������������������       �Q/?l�@B            �\@                           @��c5C @e           ��@������������������������       ��oLN��?�            �v@������������������������       ����c�@            �h@                           @��s�Z@�           �@                           �?t��P�@�           |�@                            �?F��j��	@�           p�@������������������������       ����8�	@�            �p@������������������������       �uK���	@�           �@                           �?���ܳ@`           @�@������������������������       �
f�-��@9            �Y@������������������������       �߁��F@'           ��@                           �?5|���	@�            `s@                            �? ���L�	@K            @^@������������������������       ����� 4@            �G@������������������������       �mɹ��b	@-            �R@                           !@<����@{            �g@������������������������       �-�)΃p@r             f@������������������������       ��$��� @	             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     0s@     (�@      ;@      J@     z@     @W@     ��@     �m@     H�@     �v@      ;@             �T@     �c@      @      @     �X@      "@     0}@     �D@     �q@     @T@      @              E@     �R@       @      @     �M@      �?     �Y@      >@     @Z@     �M@      @             �A@      H@       @      @      D@      �?     @X@      .@     �T@     �B@      @              "@      $@                      *@              F@      @      C@       @                      :@      C@       @      @      ;@      �?     �J@      $@     �F@      =@      @              @      :@                      3@              @      .@      6@      6@      �?               @      @                      @              @      �?      "@      @                      @      3@                      (@              @      ,@      *@      .@      �?             �D@     �T@      �?      @     �C@       @     �v@      &@     �f@      6@       @              2@      (@                      2@      @     @R@      @      H@      @                      @      @                      @              8@      �?      >@      @                      &@      "@                      ,@      @     �H@      @      2@      �?                      7@     �Q@      �?      @      5@       @     0r@      @     �`@      0@       @              "@     �D@                      (@       @     `j@      �?     @T@      $@                      ,@      >@      �?      @      "@              T@      @     �I@      @       @      6@      l@     �x@      8@     �F@     �s@      U@     �@     `h@     `�@     pq@      5@      (@     `g@     �u@      7@     �D@     �q@     �Q@     @@     �c@     @~@     �n@      (@      (@     @[@     �b@      4@      5@     �a@      E@      ^@      Y@     �a@     �a@      &@      �?      =@     �A@      @       @      E@      ,@      E@     �A@      A@      4@      @      &@      T@     �\@      0@      *@     �X@      <@     �S@     @P@     �Z@     @^@      @             �S@     @i@      @      4@     �a@      =@     �w@      M@     �u@     @Z@      �?               @      6@              $@      &@      @      *@      &@      4@      @                      S@     �f@      @      $@      `@      7@     �v@     �G@     @t@     �X@      �?      $@     �B@     �D@      �?      @      C@      *@     �G@     �B@      D@     �@@      "@      $@      .@      *@                      4@      @      (@      4@      "@      &@      @               @      @                      $@       @              "@      @      @      �?      $@      @       @                      $@      @      (@      &@       @      @      @              6@      <@      �?      @      2@      @     �A@      1@      ?@      6@      @              3@      <@      �?      @      1@      @     �A@      1@      ;@      5@      @              @                              �?      @                      @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJL�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@&��%"5@�	           ��@       	                    @�H�|�@{           6�@                           �?�����@�           Б@                           @�{���@�           �@������������������������       ��0�94@{           x�@������������������������       �F\�4Z	@r            @f@                          �1@%�z{�@�            0w@������������������������       ��mJ2@5             U@������������������������       �0$�n2@�            �q@
                           @��dAH@�           ��@                           �?<����P@�           ��@������������������������       �N����@           Py@������������������������       �e�ja-@�            v@                          �3@���L�@�            s@������������������������       �/Q,�K�@�            �i@������������������������       ���od�@C            @Y@                           @�vp�h�@;           ��@                          �<@Ej;�	@�           ��@                           �?v�En�@           ��@������������������������       �?w_s�@}             i@������������������������       ��ڱ:��@�           ��@                           �?�ڢ	�@�            �m@������������������������       �I����@,            �Q@������������������������       ��SHB�$	@l            �d@                           @��f���@�            �@                           @�{q��@           �{@������������������������       ��A���C@�            @q@������������������������       �k6[�b�@e             e@                          �:@Hۉ�2�@�             i@������������������������       �/X@\            �b@������������������������       �X0n���@%             J@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     @r@     @�@     �A@     �H@     `{@     �X@     ��@     @j@     x�@     w@      0@      @     �]@     �t@      $@      7@     �j@     �D@     8�@     @W@     @     �b@      @      @      S@     �g@      @      ,@      b@     �@@     �n@     @T@     �m@     �Z@      @      @      P@     @]@      @       @     �\@      8@     �`@     �L@     �c@     �S@      @      @     �G@     �T@      @       @      U@      (@     �Z@      C@     �a@     �P@      �?      @      1@      A@      �?      @      >@      (@      <@      3@      ,@      (@       @              (@     �Q@      �?      @      >@      "@     �[@      8@     �S@      <@                      �?      7@                      @              A@      "@      *@      �?                      &@      H@      �?      @      ;@      "@     @S@      .@     �P@      ;@                     �E@     �a@      @      "@     �Q@       @      }@      (@     Pp@     �F@      @              >@     �Z@       @              D@      @     �u@      $@     `g@      =@      �?              *@     �F@                      :@      �?      h@      "@      Y@      2@      �?              1@     �N@       @              ,@      @     �c@      �?     �U@      &@                      *@     �A@      �?      "@      ?@      @     �]@       @     �R@      0@      @               @      1@              @      8@             @U@      �?     �I@       @      @              @      2@      �?       @      @      @     �@@      �?      7@       @               @     �e@     �o@      9@      :@     �k@      M@     �q@     @]@     �s@     @k@      "@      @     @^@      e@      0@      4@     �b@      D@     �_@     �W@     @d@      c@      "@      @     �X@     �a@      ,@      &@     @^@      :@     @]@     �P@     @`@     @W@      @       @      ;@     �A@      @      �?      2@              F@      &@     �G@      $@       @       @     �Q@     �Z@      &@      $@     �Y@      :@     @R@     �K@     �T@     �T@      @       @      7@      :@       @      "@      >@      ,@      "@      <@      @@      N@      @              @      ,@              @      @              @      @      "@      7@      �?       @      0@      (@       @      @      8@      ,@      @      7@      7@     �B@       @       @      J@     �U@      "@      @      R@      2@     @c@      7@     �c@     @P@               @      6@      N@       @      @     �D@      2@     �^@      ,@      ^@     �@@               @      $@      A@               @      <@      @     �V@      @     �S@      3@                      (@      :@       @      �?      *@      (@     �@@       @     �D@      ,@                      >@      ;@      �?      @      ?@              ?@      "@      B@      @@                      0@      6@      �?              7@              <@      @      7@      <@                      ,@      @              @       @              @       @      *@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJqF�QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�9��S@�	           ��@       	                   �8@Ή�`�@g           �@                           �?��ӏ�,@�           8�@                           �?�Fkz9@C           �@������������������������       ��2�(@�            `v@������������������������       �|&�@[            �c@                           �?r�U��@�           0�@������������������������       ���Q�M	@�           ��@������������������������       ���+@w@�            �q@
                           �?,���'d	@�           H�@                          �:@ ZU�}	@<           @~@������������������������       �1R�	�e@l            �e@������������������������       �C�DM8w	@�            Ps@                            �?/E���*@O            �`@������������������������       �\��}��@            �@@������������������������       �gm��@8             Y@                           �?��_ C@D           H�@                          �2@`�I��@�           H�@                           @�P���F�?�            `p@������������������������       �����?|            @g@������������������������       �)gb*@0             S@                           �?�6�$RJ@�            0v@������������������������       ��Ű��@�            `s@������������������������       ������@            �F@                          �7@��B��@�           ��@                          �1@8kI%�\@           (�@������������������������       �aE+oI @}            `i@������������������������       ��`�:p@�           Ѓ@                           @�c�:��@�            @r@������������������������       �r�T�2�@~            �g@������������������������       ��vh�2@9            �Y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     0r@     ��@      5@      J@     �}@     @U@     Ў@      m@     Ȉ@     �u@      A@      3@     �i@     �t@      .@     �C@     �t@      Q@      v@     `f@     Pw@     @l@      ;@      (@     �^@     �n@      "@      ?@     `n@      F@      s@      Z@     �q@     �`@      *@             �E@     �S@      �?      @      L@      @     `c@      2@     �^@      <@      @              @@      Q@      �?      @      F@      @     �U@      0@     �S@      7@      @              &@      $@                      (@      @      Q@       @     �F@      @              (@     �S@     �d@       @      <@     `g@      C@     �b@     �U@     �d@     �Z@      $@      (@     �P@      [@      @      4@      b@      @@     @X@     �N@     �^@      S@      "@              *@     �M@      �?       @      E@      @      K@      9@     �D@      >@      �?      @     @U@      U@      @       @      V@      8@      H@     �R@     �U@      W@      ,@      @      R@      O@      @      @     �Q@      2@     �A@      P@      N@     �Q@      *@             �@@      ;@               @      8@      @      .@      8@      9@      (@       @      @     �C@     �A@      @      @     �G@      *@      4@      D@     �A@     �M@      @              *@      6@              @      1@      @      *@      &@      :@      5@      �?                      $@                      @      �?      @              @      @      �?              *@      (@              @      $@      @      "@      &@      3@      2@                      U@     �n@      @      *@      b@      1@     ��@     �J@     @z@      _@      @              ;@     �X@       @       @      A@      *@     0q@      3@      `@      2@                      *@      ?@               @      "@       @      d@      @      D@       @                      @      :@                      �?       @     �^@              ;@      �?                      @      @               @       @             �B@      @      *@      �?                      ,@      Q@       @              9@      &@     �\@      0@      V@      0@                      (@     �N@       @              9@      @      [@      &@     @R@      &@                       @      @                              @      @      @      .@      @                     �L@     `b@      @      &@     �[@      @     Pv@      A@     @r@     �Z@      @             �C@     �^@       @      @      N@       @     0s@      .@     �k@     �L@      @              �?      8@               @      "@             �U@      @      Q@       @                      C@     �X@       @       @     �I@       @     �k@      $@     `c@     �H@      @              2@      9@       @      @      I@       @      I@      3@     @Q@     �H@      �?              &@      2@              �?      B@             �D@      @     �I@      9@      �?              @      @       @      @      ,@       @      "@      ,@      2@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJt��vhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �5@?24�@�	           ��@       	                    �?N
���c@}           P�@                           �?��Ƚ@�           X�@                           @�� �$@�            �x@������������������������       �����@b            �c@������������������������       �<a΅n�?�            @n@                            �?\�\D��@�            �w@������������������������       �dk�Jd�@�            @i@������������������������       �	N�g�@p            @f@
                           @��8l@�           t�@                           @#M�<��@1           ��@������������������������       ���C�?@W           `�@������������������������       ����@@�            0u@                          �1@�ui@^            �c@������������������������       ��
�@            �@@������������������������       �o�Dڵ�@M            @_@                           �?���o�@B           ��@                           �?�e��;@2           �|@                          �<@h���@�            �j@������������������������       �ϯ����@q            �d@������������������������       ���^�L�@$             I@                           @�d�~@�            �n@������������������������       �eY�-@)            @Q@������������������������       ��k�8�@t             f@                          @A@� �M�'	@           T�@                           @B*�l�	@           ��@������������������������       �p_ŵ�	@�           x�@������������������������       ��!] �@           �|@������������������������       �Z��h W@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     Pr@     ��@      :@     �G@     �{@     �T@     l�@     @j@     ��@     �u@      B@      @     @]@     �s@       @      6@      j@      @@     �@     �T@     �@     �c@      1@              D@     �X@      �?      @     �G@       @     �u@      6@     �d@     �E@      @              .@      H@      �?      @      ;@       @     `g@      ,@     �Q@      8@      @              "@      1@      �?      @      .@       @      J@      *@      ?@      "@      @              @      ?@               @      (@             �`@      �?      D@      .@                      9@      I@                      4@             �d@       @     @W@      3@      �?              .@      A@                      @             @S@      @      L@      $@                      $@      0@                      *@             �U@      @     �B@      "@      �?      @     @S@      k@      @      .@     @d@      >@     0x@     �N@     �u@     �\@      *@      @      Q@     @i@      @      *@     @b@      ;@     v@      F@     �s@     �V@      @      @     �K@     �`@      @      $@     @^@      7@      p@      7@     �l@     �R@      @              *@      Q@      @      @      9@      @     @X@      5@     �U@      0@       @      @      "@      .@               @      0@      @      A@      1@      >@      7@      @               @                      �?                      *@       @      @      "@              @      @      .@              �?      0@      @      5@      .@      8@      ,@      @      "@      f@     �o@      2@      9@     `m@      I@     �s@     �_@     �q@      h@      3@              ?@     �P@       @      @      I@      @     �_@      3@     �Y@     �G@      @              6@      D@       @      @      @@      �?      @@      *@      C@      :@      @              2@      >@       @       @      =@      �?      =@      &@     �A@      @      @              @      $@              @      @              @       @      @      5@                      "@      :@                      2@      @     �W@      @     @P@      5@                      @       @                      @              <@      @      3@      @                      @      8@                      .@      @     �P@      �?      G@      .@              "@      b@     @g@      0@      3@      g@      F@     @g@      [@     @f@      b@      0@      @     `a@     �f@      (@      3@      g@      F@     @g@      [@     �e@     �a@      0@      @      Y@     @\@      "@      0@     �Z@      C@     �U@     �T@     �S@     �X@      0@             �C@     @Q@      @      @     �S@      @      Y@      :@     �W@     �E@              @      @      @      @                                              @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�c�'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?P�}� ^@�	           ��@       	                     �?�W�T��@           ��@                          �6@:��w�@�             u@                           �?�*�>@�             n@������������������������       �(f|��@2             U@������������������������       �Ty�����?c            �c@                          �<@z٭��W@=            �X@������������������������       �.�C�u&@2            @T@������������������������       ���H �@             1@
                            �?P�°�@@:           ��@                           �?�k>�Dk@�            �t@������������������������       ��/�2!F@y            @h@������������������������       �4rP���@X            �a@                          �5@�;9��S@i           �@������������������������       �y�%��4@�            0t@������������������������       �>�:H@�            �o@                           �?4-�t/@�           Τ@                           @K�*d�	@�           D�@                          �9@� ��N	@�            �n@������������������������       ���%�Z�@o            �d@������������������������       ��=��M�@0             T@                           �?�;7C�a	@@           �@������������������������       ��sO*�@�             v@������������������������       �����5	
@j           ؁@                           @P|�M�@�           X�@                           @R��B��@P           ��@������������������������       �UZ=��W@f           (�@������������������������       ����g�@�           (�@                           �?�59�FV@n            �e@������������������������       �,�����@)             L@������������������������       ���ݱ��@E             ]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     `s@     �@     �A@     �M@     `}@     @U@     �@      k@     x�@      v@      9@              X@     �e@      @      (@      ]@      "@     �z@     �I@     �p@     �U@      @              *@     �H@      �?      �?      =@              `@      ,@      R@      =@       @               @      C@                      (@             @Z@      @      H@      6@                      @       @                      @              :@      @      3@      &@                       @      >@                      @             �S@              =@      &@                      @      &@      �?      �?      1@              7@      @      8@      @       @              @      @      �?      �?      0@              7@      @      3@      @                      �?      @                      �?                       @      @      �?       @             �T@      _@      @      &@     �U@      "@     �r@     �B@     �h@      M@      �?             �C@      F@      �?       @      @@      @      V@      (@     �R@      >@      �?              8@      9@      �?      @      5@      �?     �M@      @      @@      1@                      .@      3@              �?      &@      @      =@      @     �E@      *@      �?              F@      T@       @      @     �K@      @     �j@      9@     �^@      <@                      3@      ?@                      ?@      @     `b@      $@     �Q@      $@                      9@     �H@       @      @      8@      �?     �P@      .@      J@      2@              ,@     �j@      y@      ?@     �G@      v@      S@     ��@     �d@     �@     �p@      6@      ,@      ]@     @h@      4@      5@      g@      M@      _@     �[@      e@     �a@      .@      @      >@      2@      @      @     �E@      0@      3@      4@     �K@      :@      @      @      1@      "@      @       @     �C@       @      3@      @     �A@      0@      @              *@      "@              �?      @       @              *@      4@      $@       @      $@     �U@      f@      0@      2@     �a@      E@     @Z@     �V@     �\@     @]@      "@              6@     @T@       @      @      O@      @      P@      2@      G@     �F@      �?      $@      P@     �W@      ,@      &@     �S@      B@     �D@     @R@      Q@      R@       @             �X@     �i@      &@      :@     @e@      2@     @{@      K@     �u@      _@      @             �S@      g@       @      7@     �b@      .@     px@      D@     t@     @[@       @              B@     @V@              @     @R@      *@     �b@      9@     @Z@      I@       @              E@      X@       @      0@     @S@       @     @n@      .@      k@     �M@                      4@      5@      @      @      4@      @     �F@      ,@      7@      .@      @               @      @              @      @      �?      (@      @       @      @      @              (@      0@      @              *@       @     �@@      &@      .@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ_��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �7@�ϡ��B@�	           ��@       	                    �?+NQ6�@�           ��@                          �3@Tp)���@           �@                          �1@�ߘ��@�           ��@������������������������       ��׎�)@�            �t@������������������������       �s|F�$z@�             w@                            @�9;�_�@t           (�@������������������������       �AJ΃x%@           �z@������������������������       �dk����@e            �c@
                           @�&�-@�           8�@                           �?��"p�@1           �@������������������������       ���%�sa@�            @n@������������������������       �U�u�sj@�           ��@                           @C;��i@�           X�@������������������������       �ьs��c@c            �d@������������������������       ��ȁ+�@0           @|@                           @�IT�%	@�           ܑ@                           @g�]�S�	@�           P�@                           �?,���Ӗ	@�           h�@������������������������       ���7r�	@U           x�@������������������������       ����`��@V            �_@                            �?�Mh�	@;            @W@������������������������       ����N�@             B@������������������������       ��T���T@%            �L@                          �<@r}���@�            �x@                          �9@�s[���@�             s@������������������������       ���=���@e            �d@������������������������       ���]c6@X            �a@                           �?�����O@6            �V@������������������������       ����0��@            �B@������������������������       �)C{G	@#             K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     @r@     p�@     �B@      M@     �|@     �O@     ��@     �j@     Ј@     �u@      =@      $@     @h@     �{@      4@      @@     Pr@     �A@     @�@     @\@     �@     @i@      *@      �?     �R@      k@      &@      .@      b@      7@     z@      F@      n@     �V@       @      �?      B@      Y@      @      @      R@      @      p@     �A@      b@      F@       @      �?      &@     �H@      �?      @      >@      �?      b@      0@      O@      ,@                      9@     �I@      @              E@      @     @\@      3@     �T@      >@       @              C@      ]@      @      (@     @R@      3@     �c@      "@      X@      G@      @             �@@     �V@              "@      K@      .@     �_@       @      L@      =@      @              @      :@      @      @      3@      @      @@      �?      D@      1@       @      "@      ^@      l@      "@      1@     �b@      (@     pz@     @Q@     u@      \@      @      "@     @V@      `@      @      ,@     @]@      $@     �d@      O@     �f@     @U@      @              :@      @@              �?      8@             �P@      @     @P@      6@              "@     �O@     @X@      @      *@     @W@      $@     @X@     �L@     @]@     �O@      @              ?@      X@      @      @      ?@       @     0p@      @     `c@      ;@       @              &@     �B@       @              @      �?     �Q@              A@      @                      4@     �M@      @      @      8@      �?     �g@      @     @^@      7@       @      *@     �X@     �b@      1@      :@     �d@      <@     `e@      Y@      k@     �a@      0@      &@     @R@     �[@      .@      6@     �\@      :@     @Q@     �V@     �Z@     �W@      ,@      @     �O@     @Y@      (@      6@     �X@      5@      P@     �Q@     @X@     �V@      $@      @     �K@     �S@      (@      3@      V@      .@     �D@     �N@     @R@     �Q@      "@               @      6@              @      &@      @      7@      "@      8@      3@      �?      @      $@      $@      @              .@      @      @      4@      $@      @      @               @      @      @               @      @              $@      @       @      @      @       @      @                      *@      �?      @      $@      @       @               @      9@      C@       @      @     �I@       @     �Y@      $@     �[@     �H@       @       @      0@      =@      �?      @      =@       @      V@       @     �W@      >@       @       @      &@      2@              �?      0@             �K@      �?     �C@      5@       @              @      &@      �?      @      *@       @     �@@      @      L@      "@                      "@      "@      �?              6@              ,@       @      .@      3@                      @      �?                      @              &@              @       @                       @       @      �?              3@              @       @       @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ#E�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��InD@�	           ��@       	                   �9@�%� ��@x           6�@                          �1@�o���0@0           �@                           �?��.��@�            @p@������������������������       ����
�@i            �c@������������������������       �,��违@A            �Y@                          �3@�e��@�            �@������������������������       ��ׇ�\�@           �y@������������������������       �&��E��@z           (�@
                          �:@T����	@H           ��@                           @\}x��@G            �]@������������������������       �� icg@+            �R@������������������������       ��� �3@            �F@                            �?vLs�{	@            z@������������������������       ���f@D            �[@������������������������       ���9��"	@�             s@                          �4@��7�+@0           ��@                           �?J�h�@T           �@                            @I��9��?�            �u@������������������������       ����>�G�?�            �q@������������������������       �۱����?&             M@                           @�alt�@z           P�@������������������������       �jm���@%           �}@������������������������       ��. *O�@U            �a@                          �6@�K;?�=@�           `�@                          �5@'��7I@�            `q@������������������������       �P;,=4@i            �c@������������������������       �aXj~��@G            �]@                           @��0 �@,           `}@������������������������       �2[rK�@�             r@������������������������       �
�ւk�@u            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     �@      ;@     @P@      |@      U@     8�@     `j@     ��@      w@      ?@      0@      k@     �s@      6@      I@     �r@     �I@      y@     @f@     �w@     �n@      :@      @     �b@     �o@      ,@      C@     �k@      >@     �u@      ]@     ps@      d@      5@              *@     �C@       @             �@@             �T@      &@     �L@      7@                      (@      8@       @              9@             �D@      �?      B@      1@                      �?      .@                       @             �D@      $@      5@      @              @     @a@     �j@      (@      C@     �g@      >@     pp@     @Z@     �o@     @a@      5@       @     �C@     �F@       @      @      G@      $@     �V@     �B@     �S@      K@      �?      @     �X@     @e@      $@      ?@     �a@      4@     �e@      Q@      f@      U@      4@      $@     @P@     �N@       @      (@     �T@      5@     �L@      O@      Q@      U@      @              ,@      *@       @              2@      &@      $@      6@      2@      "@       @              "@       @                      .@      &@       @      ,@      (@      @                      @      @       @              @               @       @      @      @       @      $@     �I@      H@      @      (@      P@      $@     �G@      D@      I@     �R@      @       @      @      $@       @       @      <@      @      4@      "@      *@      ,@      �?       @      H@      C@      @      $@      B@      @      ;@      ?@     �B@     �N@       @             �Q@     �l@      @      .@     `b@     �@@     ��@     �@@     �y@     @_@      @              @@     �^@       @      @      K@      @     �z@      *@      n@     �K@                       @      A@              @      ,@             �h@      @     @R@      "@                      @      @@              @      ,@              e@      @     �K@      @                      �?       @              �?                      ?@              2@      @                      8@     @V@       @       @      D@      @     �l@      $@      e@      G@                      *@     �R@                      =@      @     @f@      "@     �_@     �D@                      &@      .@       @       @      &@      @      J@      �?     �D@      @                     �C@     �Z@      @      "@     @W@      :@     �i@      4@      e@     �Q@      @              @      E@               @     �@@      &@     �X@      �?     �M@      5@      @              @      <@               @      4@       @     �E@      �?     �D@      "@      @              @      ,@                      *@      @      L@              2@      (@                     �@@     @P@      @      @      N@      .@      [@      3@     �[@     �H@      �?              8@      C@              @      B@      @     �R@      @     �P@     �@@      �?              "@      ;@      @      @      8@      $@     �@@      *@     �E@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�6!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �3@UP�\f@�	           ��@       	                    �?��n�@�           ��@                           �?0Z�H�@2           p}@                            �?�v�K@k            @e@������������������������       ��o"�@5            �U@������������������������       ��i��Y@6             U@                           @�>��p@�            �r@������������������������       �I�$��@�             j@������������������������       ��k�;N@@             W@
                           @U7��8|@_           ��@                            �?Yo�@�            �x@������������������������       �[
�>�|@F            �[@������������������������       �����\B@�            �q@                            �?[{���L@e           X�@������������������������       �"�4�S@�            �u@������������������������       ���g�� @�            �m@                           @f�kn@           :�@                           @yl��@r            �@                          �;@��	@E           Ԕ@������������������������       ��1tY�@�           ��@������������������������       �ʘbj�
@�            Pq@                            �?�q�;(@-           ؊@������������������������       ����6�@|            �h@������������������������       �Q_�O�@�           ��@                           !@pW:�	@�            �p@                          �8@10`;�;	@�            `o@������������������������       ���El@W             b@������������������������       �s����0	@A            �Z@������������������������       �ʁ�Y3@
             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@      s@     ؀@      <@      K@     p}@     �T@     ��@      m@     @�@     w@      >@      @     @R@      g@      @      .@     �_@      *@     @�@      P@     0t@     �^@      �?      @      A@     �J@       @      @     @Q@      &@     @[@      F@     �S@     �M@      �?               @      9@                      7@      @     �I@      &@     �A@      *@                      �?      *@                       @              <@      "@      2@      "@                      @      (@                      .@      @      7@       @      1@      @              @      :@      <@       @      @      G@      @      M@     �@@      F@      G@      �?       @      .@      &@       @      @      D@      @      C@      4@     �A@     �B@               @      &@      1@               @      @       @      4@      *@      "@      "@      �?             �C@     �`@       @      "@      M@       @     �y@      4@     �n@      P@                      :@     @P@              �?      :@       @     �b@      ,@     �T@      =@                       @      1@                      @              H@      @      ;@       @                      8@      H@              �?      5@       @     @Y@      $@     �K@      5@                      *@     �P@       @       @      @@             `p@      @     @d@     �A@                      @      @@       @      @      5@             �c@      �?      W@      =@                      @     �A@              �?      &@              Z@      @     �Q@      @              .@     �l@      v@      8@     �C@     �u@     @Q@     �|@      e@     P~@     �n@      =@      (@      i@     �s@      5@      C@     �r@      K@      z@     ``@      }@      l@      .@      &@     �c@     �h@      *@      @@      j@      C@      f@     �[@     @k@     �c@      .@      @      `@      c@      @      5@      f@      8@     �b@      V@     �f@      [@      *@      @      >@      F@      @      &@      ?@      ,@      <@      6@     �A@      H@       @      �?      E@     @]@       @      @     �V@      0@      n@      5@      o@      Q@                      *@      1@       @              <@       @     �N@      @      I@      1@              �?      =@      Y@      @      @     �O@      ,@     �f@      ,@     �h@     �I@              @      ?@      D@      @      �?     �F@      .@     �C@     �B@      3@      6@      ,@      @      ;@     �C@      @      �?     �E@      &@     �C@      B@      3@      5@      "@              $@     �@@              �?      @@      @      7@      (@      $@      *@      @      @      1@      @      @              &@      @      0@      8@      "@       @      @              @      �?                       @      @              �?              �?      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ}rfOhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��:�9@�	           ��@       	                    �?��jX<	@�           �@                           �?�ia\�@p           ��@                            @/�����@p            �d@������������������������       �zu�^<�@S             `@������������������������       �ڼoc�@            �B@                           @�@���@            �x@������������������������       �[<�$�!	@;            �V@������������������������       ���(�Y�@�            s@
                           @�`T�	@c           ��@                          �9@����		@h            �@������������������������       ���Vn@            z@������������������������       ��\�Զ@g             d@                           @����_'
@�            y@������������������������       ��s%���	@�            �w@������������������������       �Ϝ��@             3@                          �5@�sw�W@�           ��@                           @-��5s@�           �@                            �?�]�:@|            �@������������������������       ����ނ@n            �g@������������������������       ��3 4x@           Pz@                            �?T���~�@!           �@������������������������       ��
�$Q��?v             g@������������������������       �d};ə@�           H�@                           �?AR�*��@0           �@                          �=@� ��и@�            �m@������������������������       �J\v��(@�            �j@������������������������       �P:&У@             8@                           @� j9��@�           ��@������������������������       �b� �9@�           p�@������������������������       �I5�b�@             C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     8�@      ?@      I@     �{@     �S@     `�@     @k@      �@     v@      B@      *@     �d@     �n@      6@      :@     �k@      I@     �j@      _@     �o@     �e@      ;@       @      D@     @W@      @      @      V@      $@     �Z@      D@     @Z@     �N@      @              ,@      =@                      8@              D@      @     �G@      "@                      *@      3@                      5@              ?@      �?     �A@      "@                      �?      $@                      @              "@       @      (@                       @      :@      P@      @      @      P@      $@     �P@     �B@      M@      J@      @       @      @      @      @      �?      0@      @      "@      "@      7@      $@       @              5@     �L@       @      @      H@      @     �L@      <@     �A@      E@      @      &@     �_@     @c@      1@      3@     �`@      D@      [@      U@     �b@     @\@      6@      @      Q@     @X@      $@      (@     �T@      5@     �S@      =@     @Y@      P@       @      �?      L@     �K@      "@      $@     @Q@       @     �P@      2@     @T@      C@      @      @      (@      E@      �?       @      ,@      *@      *@      &@      4@      :@      @      @      M@     �L@      @      @      J@      3@      =@     �K@     �G@     �H@      ,@      @      L@     �L@      @      @      H@      3@      =@      K@     �F@      G@      &@      @       @                              @                      �?       @      @      @       @     ``@      s@      "@      8@     �k@      =@     ��@     �W@     8�@     `f@      "@             �F@     �i@      @      0@      \@       @     ؁@      F@     `w@     @W@      @              9@      Y@      �?      @      N@      @     �h@      @@      `@     �J@      �?              @      9@                      (@      @     @Q@      $@      G@      7@                      6@     �R@      �?      @      H@      @     @`@      6@     �T@      >@      �?              4@      Z@      @      &@      J@      �?     @w@      (@     �n@      D@      @              �?      .@                      &@              [@       @     �D@      @                      3@     @V@      @      &@     �D@      �?     �p@      $@     �i@      A@      @       @     �U@      Y@      @       @      [@      5@     `k@      I@      j@     �U@      @              0@      9@                      (@      @     �T@      @     @R@      ,@      @              .@      8@                       @      @      T@       @      Q@      &@                      �?      �?                      @      �?       @      @      @      @      @       @     �Q@     �R@      @       @      X@      .@      a@      F@      a@      R@      �?       @      M@     �R@       @       @     �V@      *@      a@      B@     @`@      R@      �?              (@      �?       @              @       @      �?       @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@>����b@�	           ��@       	                     @x�>�@P           ��@                          �1@d�N��@�           ��@                           �?3 �$U@           {@������������������������       �2bN��?q             f@������������������������       �4�u?��@�             p@                          �4@�m���@�           ��@������������������������       �4���@5            �@������������������������       �l ��?�@�            �o@
                           �?� �f�5@b           @�@                           �?��2���@y            �g@������������������������       ����0�g�?             B@������������������������       ���<�B@a             c@                           �?f.l�Ex@�            �v@������������������������       �w�q�8	@�            @l@������������������������       ��Y{���@S             a@                           �?������@l           ě@                          �<@��w	@1           8�@                           �?�U��>:	@�           ��@������������������������       ��we�$@z            �f@������������������������       ��G@"�	@7           �}@                           �?�Ϫ�5�@�            `j@������������������������       ��qqh.�	@/             S@������������������������       �d���M@Q            �`@                           @�9/�Z@;           P�@                          �7@=:'��@�           X�@������������������������       ����!�@�            `q@������������������������       �/�6d��@?           P@                          �:@u9r)U0@G            �_@������������������������       �Lf�!�g@1            �V@������������������������       � �'�j�@            �B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        &@     @r@     �@     �C@     �K@     �|@     @W@     x�@     �k@     8�@     �w@      ?@      @     �Z@      r@      .@      5@     @j@      A@     `�@     �X@     �~@      e@      .@             �Q@     �j@      $@      (@     �c@      9@      �@     �Q@     `v@      \@      "@              "@      M@              @     �B@      @      g@      &@      Z@      6@      �?              @      3@               @      0@             �X@              ?@      @      �?              @     �C@               @      5@      @     �U@      &@     @R@      0@                      O@     `c@      $@       @     �]@      6@     �v@     �M@     �o@     �V@       @             �I@     �\@      "@      @     �V@      $@      s@      J@     �f@     �Q@       @              &@     �D@      �?      @      =@      (@      N@      @     �Q@      4@              @     �A@     �R@      @      "@      K@      "@      a@      =@     �`@      L@      @              (@      1@               @      @       @     �U@      @      H@      (@                               @                                      1@      �?      $@                              (@      "@               @      @       @     @Q@       @      C@      (@              @      7@      M@      @      @     �G@      @      I@      :@     �U@      F@      @      @      4@      ;@      @      @      C@      @      7@      0@     �I@      =@      @              @      ?@      �?      @      "@              ;@      $@     �A@      .@      @      @     @g@     @l@      8@      A@     �o@     �M@     0t@     �^@     �s@     �j@      0@      @     �X@     �^@      0@      6@     �`@      @@     �Y@     @S@      ]@     �`@      &@       @     @T@     �X@      (@      ,@     �Y@      4@      V@      J@     @Y@     �S@      &@      �?      :@      <@       @      @      8@              A@      $@      D@      ,@      �?      �?     �K@     �Q@      $@      &@     �S@      4@      K@      E@     �N@     @P@      $@      @      2@      8@      @       @      ?@      (@      .@      9@      .@      L@               @      @      *@      @      @      (@      @       @      @      @      *@              �?      *@      &@      �?      @      3@      @      @      3@      &@     �E@               @     �U@      Z@       @      (@     �]@      ;@     �k@      G@     �h@     @S@      @       @     �O@     �U@      @      (@     �Z@      5@      h@     �A@      g@     �Q@       @              ?@     �@@      @      @      <@      @      X@      @     �I@      4@       @       @      @@      K@               @     �S@      1@      X@      ?@     �`@      I@                      8@      1@      @              *@      @      <@      &@      .@      @      @              (@      0@      @              @      @      ;@      $@      @      @      @              (@      �?                       @      �?      �?      �?      $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�>�zhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��Q�E@�	           ��@       	                    �?�h��@�           t�@                           �?M\{A�[@,           `}@                            @d��T�f@p            �g@������������������������       ���j�@N            �a@������������������������       ��:#>�@"            �I@                            �?XRj���@�            pq@������������������������       ����5;@9             U@������������������������       �f�%�@�            `h@
                           �?fѧY�e@�           8�@                            �?0(���@           py@������������������������       ��/B���?>             X@������������������������       �>q�@@�            ps@                          �=@{�fy.@�             s@������������������������       ��7"u�r@�            0r@������������������������       ��g�L@
             *@                          �1@L�:��@�           X�@                           @��/�B@�            �v@                          �0@+��3@$             K@������������������������       �f�#G 5�?             *@������������������������       �:p��@            �D@                           @��p�^@�            `s@������������������������       �V,�@y            �g@������������������������       ���}�_@O            �^@                          �;@�
�}�y@�           ��@                           @Jm��n%@�           ��@������������������������       ���ɦrB	@�           ��@������������������������       ���籝@           ��@                           �?��;=k	@�            �u@������������������������       �2�����	@v             g@������������������������       ��i~.@]            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@      s@     ��@      ;@      H@     �|@     @T@     Ȏ@     @k@      �@     `w@      9@       @      U@     �d@       @      @     �Z@      $@     `y@     �D@     �q@     �Q@      @       @     �G@      V@              @      M@      �?     �U@      <@     �[@     �F@       @       @      4@      @@                      9@              E@      @     �H@      .@      �?       @      1@      3@                      7@              9@      @     �A@      ,@      �?              @      *@                       @              1@      �?      ,@      �?                      ;@      L@              @     �@@      �?      F@      7@     �N@      >@      �?              @      3@              �?       @      �?      ,@      @      9@      @                      4@     �B@               @      9@              >@      4@      B@      8@      �?             �B@     �S@       @      @      H@      "@      t@      *@     `e@      :@      @              5@      J@              @      B@      @     �h@      @      R@      *@                              @               @      $@       @     �L@              (@      @                      5@     �F@              �?      :@      @     �a@      @      N@      @                      0@      ;@       @              (@      @     �^@      @     �X@      *@      @              0@      ;@       @              $@      @     �]@      @     �X@      &@      �?                                               @              @      @      �?       @       @      7@     �k@     �v@      9@      E@     0v@     �Q@     �@      f@     X�@     �r@      4@              1@     �K@       @       @      @@      �?     �_@      1@     �U@      :@                      @      @                      �?              6@      @      "@      @                       @      �?                      �?               @                      �?                      @      @                                      ,@      @      "@      @                      &@     �H@       @       @      ?@      �?      Z@      &@     @S@      6@                      @      <@       @      �?      9@              N@              K@      (@                      @      5@              �?      @      �?      F@      &@      7@      $@              7@     `i@     0s@      7@      D@     0t@     �Q@     P|@      d@     P}@     Pq@      4@      *@     �d@      p@      1@      ?@     pq@      L@     z@     �a@     �y@     �j@      2@      &@     @]@     �d@      (@      ;@     `i@     �F@      d@     @\@     �g@      b@      .@       @     �G@     �W@      @      @      S@      &@     p@      =@     �k@      Q@      @      $@     �C@     �H@      @      "@      F@      ,@      B@      2@     �L@     @P@       @      $@      2@      8@      @      @      ,@      $@      1@      ,@      4@      G@       @              5@      9@      �?      @      >@      @      3@      @     �B@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ@�{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��LS�P@�	           ��@       	                    @xZy@=           l�@                           �?�;_Ȯ@�           �@                           �?���+4@�            �t@������������������������       �+�nE`C@�            �k@������������������������       ���E��@E            �[@                           �?��d��R@�           `�@������������������������       �=_gs@�            Pp@������������������������       �Ê��~5@4           p~@
                          �4@�ôQ�@�           �@                          �0@<wO�
@4           h�@������������������������       ��p��%��??            �Y@������������������������       ����.y@�           0�@                            �?{��}�@b             b@������������������������       �p��^+�?            �B@������������������������       ����@L            �Z@                          �<@$/Mԣ�@j           L�@                           �?��h@�           ��@                           �?���g�	@�           h�@������������������������       �E9�@�            p@������������������������       �=����	@           �|@                            �?��tZp;@�           ��@������������������������       ���N��6@�            Px@������������������������       �Հ@�            �v@                           @	��a6	@�            Pu@                            �?�O$�p@�            �p@������������������������       ��L*=�@W            �`@������������������������       ���!@U            �`@                           @2�Ǟ�	@5            @S@������������������������       �����Λ	@%            �L@������������������������       �Se���?             4@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     `s@     h�@      9@     �I@     }@     �S@     �@     �k@      �@     pv@      A@      @     �\@     Ps@      @      7@     �l@      :@     `�@     @U@     @z@     `c@      *@      @     �U@     `d@      @      .@      e@      3@     @n@     @S@     @g@     @Z@      $@              ?@     �C@               @     �A@      @     @Z@      0@     @R@      =@                      ,@      ;@               @      3@       @     �P@      (@     �J@      ;@                      1@      (@                      0@      �?     �C@      @      4@       @              @     �K@      _@      @      *@     �`@      0@      a@     �N@     @\@      S@      $@      @      1@     �M@       @       @      P@       @     �B@      4@      5@      :@      �?      �?      C@     @P@      @      &@     @Q@       @      Y@     �D@      W@      I@      "@              <@     @b@       @       @     �N@      @     �}@       @     @m@      I@      @              ;@      _@       @       @     �G@             `z@       @     `h@      F@                      �?      3@                      �?             �P@              (@      @                      :@     @Z@       @       @      G@             @v@       @     �f@      D@                      �?      6@                      ,@      @      J@             �C@      @      @                      @                      "@              1@              @                              �?      2@                      @      @     �A@              @@      @      @      ,@     �h@     �q@      2@      <@     �m@      J@     Ps@      a@     �s@     �i@      5@      "@     `c@     `k@      *@      4@      h@      D@     pq@     �[@     Pq@     @a@      1@      "@     �W@     �\@       @      2@     �Z@      ;@      R@     �Q@     @\@     @Q@      ,@      �?      :@     �E@      �?      @     �F@      @      A@      1@      G@      9@       @       @      Q@      R@      @      &@      O@      7@      C@      K@     �P@      F@      @             �N@      Z@      @       @     @U@      *@     �i@      D@     �d@     @Q@      @              @@     �F@      @       @     �D@      "@     �\@      6@     @V@      =@       @              =@     �M@       @              F@      @      W@      2@     �R@      D@      �?      @     �D@     �N@      @       @      F@      (@      >@      :@     �C@     �P@      @      �?      9@      K@      @      @      B@       @      5@      2@      >@     �L@       @               @      7@              @      "@      @       @      $@      4@     �E@       @      �?      1@      ?@      @      @      ;@       @      *@       @      $@      ,@              @      0@      @              �?       @      @      "@       @      "@      "@       @      @      $@      @              �?      @      @       @       @       @      "@       @              @      �?                      @              �?              @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�_��^@�	           ��@       	                     @���E�@           ��@                           @�[6ș�@@           ��@                          �<@��A�@           0|@������������������������       �f�[o��@�            @y@������������������������       �o5���	@            �G@                          �5@��,o�@.           P}@������������������������       �J�*L�X�?�            �t@������������������������       ���Erx�@W            �`@
                           �?-8K�ǭ@�            �t@                          �7@��2գ�@|             h@������������������������       �l��T��@U            �_@������������������������       ��P6[��@'            �P@                          �:@Ȍ[t%�?X            @a@������������������������       ���8��]�?P            �_@������������������������       � ۉ����?             &@                           @ǻT71@�           ̤@                          �2@�?�(Y	@�           ��@                           �?��zeA�@�            0s@������������������������       ����A"@�            @h@������������������������       �&�v7�~@E            @\@                            �?:\aR�	@           ��@������������������������       �cBЋ�	@�           ؄@������������������������       ��Z�?#	@w           ��@                           @���T�"@�           �@                           �?ee�7��@�           �@������������������������       ���#�@?            }@������������������������       ��:h�Q@A            @                            �?��:z�@R            ``@������������������������       ����&@+            �Q@������������������������       ��uJ�=�@'             N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     ps@     �@      ;@      J@     }@     @T@      �@      i@     ��@     Px@      =@      �?     �S@      f@      @      1@     @W@      ,@     �{@     �H@     0r@     �S@       @      �?     �H@      `@      �?      (@     �P@      *@     @t@      A@     `l@      O@       @      �?     �A@      P@              &@      F@      @     �Z@      7@     �\@     �F@       @      �?      >@      M@              &@     �D@      @     @Z@      .@     �[@      :@      �?              @      @                      @               @       @      @      3@      �?              ,@      P@      �?      �?      7@       @      k@      &@     @\@      1@                      $@     �A@              �?      ,@             �g@      @      R@      "@                      @      =@      �?              "@       @      =@      @     �D@       @                      =@     �H@      @      @      :@      �?     �^@      .@      P@      0@                      9@     �C@      @      @      2@      �?      K@      (@      8@      (@                      0@      :@              �?      @      �?     �E@      @      4@      @                      "@      *@      @      @      (@              &@      @      @      @                      @      $@                       @             @Q@      @      D@      @                      @      $@                      @              P@      �?      D@      @                      �?                              @              @       @                              8@      m@      w@      7@     �A@     @w@     �P@     (�@      c@     ��@     ps@      ;@      8@     @e@     �l@      0@      <@     @n@      M@     �h@     �_@      o@      j@      5@      @      >@      I@               @     �F@      @     �Q@      9@     �I@      ;@              @      8@      >@              �?     �C@       @      6@      *@      C@      6@                      @      4@              �?      @      �?     �H@      (@      *@      @              5@     �a@     @f@      0@      :@     �h@     �K@     �_@     �Y@     �h@     �f@      5@      "@     �Q@     �U@      @      6@     @W@      @@     �O@     �Q@      [@     �W@      &@      (@     @Q@      W@      "@      @      Z@      7@     �O@      ?@     �V@      V@      $@             �O@     �a@      @      @     @`@      "@      t@      9@     �q@     �Y@      @             �I@      `@      @      @      [@      @     r@      7@     Pp@     �T@      �?              =@     �M@       @      @     @P@      �?     ``@      @     �^@     �E@      �?              6@     @Q@      @      �?     �E@      @     �c@      0@     @a@     �C@                      (@      (@      �?      �?      6@       @      ?@       @      7@      4@      @              @      @              �?      @       @      6@       @      &@      1@                      @       @      �?              1@              "@              (@      @      @�t�bub�~     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJH<QhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @h6;� @�	           ��@       	                    �?̀6�F�@x           j�@                          �:@q!�<	@            |�@                            �?	�Y��@;           ��@������������������������       �����@�            �x@������������������������       ��;��@A           ��@                           �?�ӌ~��	@�            �s@������������������������       �n�<<�@3             U@������������������������       ��4�i�Z
@�            �l@
                            @_Wȧi8@x           ��@                          �=@R+{�8@           �{@������������������������       �� s��@           z@������������������������       ��wg=��@             :@                           �?��%$i�@h            `c@������������������������       ��E,�TF@%             K@������������������������       �@�23ͩ@C            @Y@                          �6@
�h��@           P�@                           @�l�� )@�           �@                           @�1P�@�           ܑ@������������������������       ��ڛ(�@�           8�@������������������������       ��WH�@7            @������������������������       �+�%W�@
             0@                            @3|���@@           h�@                           @�*�v�@�            �y@������������������������       �9N"��@�            �x@������������������������       ��ڇ8�E@             (@                           @0�\��@A            �\@������������������������       �7�?�@             G@������������������������       �n�%��@&            @Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@     0r@     �@      @@      G@     �{@     �V@     <�@      h@     ��@     �t@     �@@      3@      j@     0v@      =@      B@     �r@     @S@     Py@     �c@     �x@     �j@      ?@      3@     �d@      q@      :@      <@      m@      L@     �o@      ]@      q@     �d@      ;@      "@      `@     �m@      .@      9@      h@      C@      k@     �V@     �m@     �Y@      9@             �J@      L@      @      @     �L@      @      S@      @@     �S@      1@      $@      "@      S@     �f@      &@      4@     �`@      ?@     �a@      M@      d@     @U@      .@      $@      B@     �@@      &@      @      D@      2@      B@      :@      A@     �O@       @      �?      @      "@              �?      .@       @      .@       @      (@      5@              "@      >@      8@      &@       @      9@      0@      5@      8@      6@      E@       @              F@     �T@      @       @     @Q@      5@      c@      D@     @_@     �H@      @             �B@     �J@      �?      @     �L@      2@     @[@      =@     @X@     �@@      @             �A@     �J@      �?      @      K@      $@     �Z@      7@     �W@     �@@       @               @                      �?      @       @       @      @       @               @              @      >@       @      @      (@      @     �E@      &@      <@      0@                       @      *@       @              @      @      (@      @      (@      @                      @      1@              @      "@              ?@       @      0@      (@                     �T@     �k@      @      $@     @b@      ,@     Ѓ@      B@     0z@     �\@       @             �C@     `e@       @      @     @U@      @     �~@      .@     @q@     �P@       @             �C@     @e@       @       @      T@       @     �~@      .@      q@      P@       @              <@     �U@       @             �C@       @      s@      (@      b@      ;@      �?              &@     �T@               @     �D@             �g@      @     �_@     �B@      �?                      �?              �?      @      @                      @       @                     �E@      J@      �?      @     �N@      "@     `a@      5@     �a@     �H@                     �B@      I@              @     �H@      @     �W@      (@     �\@      D@                      @@      I@              @      H@      @     @W@      $@     @\@      D@                      @                              �?      �?       @       @      �?                              @       @      �?      �?      (@       @      F@      "@      =@      "@                       @      �?                      �?       @      2@      "@      *@                              @      �?      �?      �?      &@              :@              0@      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��r<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���uRn@�	           ��@       	                     �?���@B           ��@                           �? �U��@           �z@                           �?B����@r            @e@������������������������       ���f �a@4            �S@������������������������       �-0):@>             W@                          �<@�շ�@�            Pp@������������������������       ��^^Nc�@�            �n@������������������������       ��bN�� @	             ,@
                           @�rL��@/           ��@                           �?�p1��
@"           H�@������������������������       ��@w�%	@�            �p@������������������������       ��� ��@s            �@                           @v౛N+@           @y@������������������������       ��͛Vm@]            @b@������������������������       ��m�ߺt@�             p@                           �?�N�{�@�           :�@                            �?% ���@{           0�@                          �2@��SsҒ@x            �h@������������������������       �B=g�;#�?'            �Q@������������������������       �Ӗ�_�#@Q            �_@                           @qZ��`@            z@������������������������       ��m���[@�            �i@������������������������       �����c%�?w            �j@                          �3@�:��@           ܘ@                          �1@9>�=g:@=           0~@������������������������       ��F�-)@�             h@������������������������       �B�;L�@�             r@                           @�����@�           P�@������������������������       ���W�N�@�           x�@������������������������       �'�=�vM@             K@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     ��@      :@     @R@     �|@      Y@     ��@      l@     `�@     �w@      7@      @      `@     �l@      &@      B@     `i@      B@     @     @Q@     �s@     `d@      (@      @      ;@      P@              @     �J@       @     �^@      @@     @V@      8@      @      @      3@      =@              �?      :@       @      8@      :@      5@      "@      @      @      @      "@                      6@      @      0@       @      @       @       @              .@      4@              �?      @      @       @      2@      ,@      @      �?               @     �A@              @      ;@             �X@      @      Q@      .@                      @      =@              @      8@             �X@      @     �P@      *@                      �?      @                      @                               @       @              @     @Y@     �d@      &@      ?@     �b@      <@     pw@     �B@     �l@     `a@      "@      @      M@     �\@      $@      ,@     @V@      5@     �q@      1@     �e@     @V@      �?      @      9@     �@@      @       @      D@      .@     �H@      &@      A@     �D@      �?             �@@     �T@      @      @     �H@      @     @m@      @     `a@      H@                     �E@     �H@      �?      1@     �N@      @      W@      4@      L@      I@       @              &@      1@              @      9@      @      7@      @      >@      1@      @              @@      @@      �?      &@      B@      @     @Q@      *@      :@     �@@      �?      @      e@     �r@      .@     �B@     �o@      P@      �@     `c@     �|@     @k@      &@              D@     @V@      @      �?      H@      @     �j@      1@     `c@      E@      �?              .@      :@      @              .@      @      R@      @     �D@      0@                      @      @                       @              G@              @      @                      $@      4@      @              *@      @      :@      @      B@      $@                      9@     �O@              �?     �@@             �a@      (@     �\@      :@      �?              5@      B@              �?      =@              E@       @      I@      2@                      @      ;@                      @             @Y@      @      P@       @      �?      @      `@     �j@      (@      B@     �i@     �N@     �r@     @a@     0s@      f@      $@       @      8@     �P@      @       @      :@       @      b@      @@      [@      N@       @              "@      <@              �?       @             �Q@       @      I@      3@               @      .@      C@      @      @      2@       @     �R@      8@      M@     �D@       @      @     @Z@     `b@      "@      <@     `f@     �J@      c@     �Z@     �h@      ]@       @      @      W@     �a@      @      <@     �d@      I@     �b@     �X@      h@      ]@       @      �?      *@      @      @              ,@      @       @      @      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ1�_OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��`Z�c@�	           ��@       	                   �3@�w�@A           ��@                            �?�p�bZ�@�           ��@                          �1@g=�ɿ@b            �c@������������������������       ��OƼ�@.            �S@������������������������       ��)~lP@4            @S@                            @�T�*s�@3            ~@������������������������       ���8")@�            �t@������������������������       �Qi��'@l            @c@
                           @e���\@�           �@                           �?�\���z	@�           X�@������������������������       �/=7��@�            @m@������������������������       ����aF�	@*           ~@                           @<���F�@�            `w@������������������������       ���Z^@�            @q@������������������������       ��@y7��@:            �X@                           �?J���`�@d           �@                            �?w1e���@d           �@                          �7@
�\޺b@�             r@������������������������       ��n$Q��@�            �k@������������������������       �ʭ�B@0            �P@                            @��%�V@�             p@������������������������       ��*i6@@            @X@������������������������       �[x��ё@b            �c@                           �?�	���z@            ��@                           @Sڧ�@G             ^@������������������������       �y��k�@@            �Y@������������������������       �F���D�?             1@                            �?�(��D@�           ��@������������������������       ������@�           ��@������������������������       ��C���s@�           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     0q@     ��@      A@      N@     `z@     �U@     X�@     `k@     ��@     `w@     �C@      @      \@     Pq@      .@      7@      h@     �A@     p~@      V@     `t@     �b@      0@      �?      9@      W@      �?      @     �J@      @     Pp@      8@     @`@      E@      �?               @      0@                      2@       @     @P@       @     �B@      @      �?              �?      @                      *@       @      C@      �?      (@      @                      �?      "@                      @              ;@      @      9@       @      �?      �?      7@      S@      �?      @     �A@       @     �h@      0@     @W@     �A@                      1@     �H@      �?      @      :@             �a@      "@     �M@      5@              �?      @      ;@                      "@       @      K@      @      A@      ,@              @     �U@      g@      ,@      3@     `a@      ?@     @l@      P@     �h@     �Z@      .@      @     @Q@     �\@      &@      1@     �Y@      :@     �\@     �K@     �Z@     @S@      .@      �?      0@      6@       @      @      ?@      �?     �S@      .@      G@      0@      �?      @     �J@     @W@      "@      (@      R@      9@     �B@      D@      N@     �N@      ,@              2@     �Q@      @       @      B@      @     �[@      "@     �V@      >@                      (@      K@               @      9@       @     �X@      @      P@      *@                      @      0@      @              &@      @      *@      @      :@      1@              "@     `d@     �q@      3@     �B@     �l@      J@      �@     ``@     �~@      l@      7@              F@      R@               @      E@      �?      h@      $@      b@      A@      @              3@      H@               @      1@      �?      X@      @     @U@      .@       @              .@      >@                      (@             �U@      @     �P@       @                      @      2@               @      @      �?      "@      �?      2@      @       @              9@      8@                      9@             @X@      @      N@      3@      �?              *@       @                      *@              @@      �?      5@       @      �?              (@      0@                      (@             @P@      @     �C@      &@              "@     �]@     �j@      3@     �A@     �g@     �I@     0t@     @^@     �u@     �g@      4@      �?      1@      @              "@      3@      @       @      1@      7@      ,@              �?      *@      @              "@      0@      @       @      *@      7@       @                      @                              @                      @              @               @     �Y@      j@      3@      :@      e@      G@     �s@      Z@     `t@      f@      4@       @     �L@     �Y@      (@      0@     �S@      5@     �c@      K@     �g@     �Y@      @      @     �F@     @Z@      @      $@     �V@      9@     �c@      I@      a@     �R@      ,@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJY�lvhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��ȟ�H@�	           ��@       	                    @��"Q�@q           �@                           �?)����@�           ��@                           �?�1.�h@�           �@������������������������       ���Yy�@�            �m@������������������������       ��r+�Do@4           @}@                           �?����y�@�            0v@������������������������       �л �Q�@Z            �b@������������������������       ���`jO@�            �i@
                           �?e	�\@�           t�@                           @"T�O��?           `z@������������������������       �������?�            @r@������������������������       �RrI@S            @`@                           @�']��w@�           ��@������������������������       �����"�@l            `f@������������������������       ��5�M@W            �@                           �?��lH�@R            �@                           �?�@k~�	@           x�@                          �9@?�OK�k@�            pp@������������������������       �z�^#�@d            @c@������������������������       �G�~qJ@N            @[@                           @`H��\ 
@i           @�@������������������������       ��O9#��	@G           ��@������������������������       �I0"�@"             I@                          �<@�� |��@7           ȋ@                           �?�H���
@�           ��@������������������������       �&���D@�            �u@������������������������       �cz)L=@�            �y@                           �?Pl�5�@T            ``@������������������������       ���/��P@            �F@������������������������       �;f��@7            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      t@     @�@      A@      F@     @{@     �T@     Џ@     @j@     ��@     �u@      A@       @     @^@     u@      1@       @      j@      ;@     Ѕ@      X@     �~@     @c@      *@       @     �P@     `e@      *@      @     �a@      3@      k@     �S@     `l@      Y@      "@       @      K@     �Y@      $@      @      [@      (@     @]@     �I@     �c@      R@      "@              3@     �D@       @      �?      7@      @      M@      1@      K@      1@       @       @     �A@     �N@       @      @     @U@      "@     �M@      A@      Z@     �K@      @              *@     @Q@      @      @     �A@      @      Y@      <@     @Q@      <@                      @      @@                      5@      @      E@      &@      2@      *@                      @     �B@      @      @      ,@      �?      M@      1@     �I@      .@                      K@     �d@      @      �?     @P@       @     ~@      1@     pp@      K@      @              1@     �Q@                      1@      �?     �m@      @      O@      (@       @              $@     �E@                      ,@      �?      f@      �?      C@       @                      @      ;@                      @              N@      @      8@      @       @             �B@      X@      @      �?      H@      @     �n@      *@      i@      E@       @              ,@     �@@                      3@      @      L@      @      @@      (@       @              7@     �O@      @      �?      =@       @     �g@      @      e@      >@              &@     �h@     �n@      1@      B@     �l@      L@      t@     �\@     �r@     �g@      5@      &@     @_@     �_@      *@      6@     @]@     �C@     �V@     @R@     �X@     �\@      2@      @      9@      C@      �?      @     �A@      "@     �H@      *@      D@     �E@       @              5@      7@      �?      @      8@      �?      C@       @      6@      1@      �?      @      @      .@              �?      &@       @      &@      &@      2@      :@      �?       @      Y@      V@      (@      1@     �T@      >@     �D@      N@     �M@     �Q@      0@      @     �W@     @T@      (@      1@     @S@      =@      B@     �H@      L@     @Q@      "@      @      @      @                      @      �?      @      &@      @       @      @             �R@     @^@      @      ,@     �[@      1@     �l@     �D@     �h@     @S@      @              M@      \@      @      "@      T@      &@     @j@      A@     @f@      N@       @              9@      I@              @     �F@             @Z@      2@     �S@      4@       @             �@@      O@      @      @     �A@      &@     @Z@      0@     �X@      D@                      0@      "@              @      ?@      @      4@      @      3@      1@      �?               @      �?              @      @      @       @      @      *@       @      �?              ,@       @                      9@      @      (@      @      @      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ[�1
hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�{��R@�	           ��@       	                   �2@�o4,J@           ̒@                          �1@H� ~B@           �y@                           @l80a2v�?�            �n@������������������������       �!�����?�            �i@������������������������       ������@             D@                           @��$��@a            �d@������������������������       �s6��1�@0             T@������������������������       ��G�����?1            �U@
                          �>@b�u�*i@           ��@                          �3@R��K�@�           (�@������������������������       �;�QH�@P            @_@������������������������       �=4���U@�           @�@                          @@@؟���_@             I@������������������������       ���E@             ?@������������������������       ���D٢U @             3@                           �?x�J@�           ,�@                          �:@�	�}�	@�            �@                            �?X1$�	@3           (�@������������������������       ��T�&x�	@�            pq@������������������������       ��O���5	@�           p�@                           @sU�>�^
@�            0p@������������������������       ���{��	@!             I@������������������������       ����r	@y             j@                           @K��u{
@�           8�@                           @����e�@b           0�@������������������������       ��A���b@�           ��@������������������������       �s����@�           h�@                            �?w]Ye��@x            @h@������������������������       ��A�1g�@             H@������������������������       �]���U�@[            @b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@      @@      O@     @{@     �V@     ��@     @k@     0�@     �u@      ;@      �?     �P@     �b@      �?      $@     �[@      *@      |@     �F@     �q@     �R@      @              @     �G@              @      D@              j@       @      S@      5@      �?              @      ;@                      5@             �a@      @     �C@      @      �?              @      7@                      (@             �_@      @     �@@      @                              @                      "@              .@       @      @      @      �?              @      4@              @      3@             �P@      @     �B@      ,@                      @      *@              @      3@              *@      @      .@      $@                              @                                      K@              6@      @              �?      N@     �Y@      �?      @     �Q@      *@     �m@     �B@     �i@      K@       @      �?      L@     �X@      �?      @     �M@      *@     @m@      =@     @h@      G@       @              &@      &@                      @      �?     �@@      @     �H@      &@              �?     �F@      V@      �?      @      K@      (@      i@      9@      b@     �A@       @              @      @                      (@              @       @      $@       @                      @                              @              @      @      @      @                              @                      @                      �?      @       @              3@     �l@     �w@      ?@      J@     Pt@     @S@     ��@     �e@     p�@     q@      8@      3@     �a@     �b@      3@      ;@     �c@      J@     �`@     �Z@     `g@      b@      5@      @     �^@     @]@      (@      7@      `@     �A@     �Z@     �R@      d@     @X@      2@      @     �F@      =@       @      &@     �B@      @     �D@      @@      E@      7@      "@      @     @S@      V@      $@      (@      W@      >@     @P@     �E@     �]@     �R@      "@      *@      4@     �@@      @      @      >@      1@      :@      @@      :@      H@      @      @      @       @      �?      �?      @      @      �?      @      &@      @      @      "@      *@      ?@      @      @      ;@      (@      9@      9@      .@     �E@                     @V@      m@      (@      9@     �d@      9@      {@     �P@     0w@      `@      @             @P@     �i@      "@      6@     `a@      5@     �w@     �I@     �u@     @\@       @             �@@      X@               @     �R@      3@     �c@     �@@     �`@      I@       @              @@     �[@      "@      ,@      P@       @      l@      2@     �j@     �O@                      8@      ;@      @      @      ;@      @     �H@      .@      :@      .@      �?              @      @      �?      @               @      "@      $@       @      $@                      2@      6@       @              ;@       @      D@      @      8@      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJR�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��߉�b@�	           ��@       	                   �1@ky�}Ѭ@[           ��@                           @�?ލ˽@�           ��@                           �?�S�G�@�             o@������������������������       ��7d[��@A            @X@������������������������       ��!H�@e             c@                           @�J�6��?�            �u@������������������������       �Ǘ �@��?�            pp@������������������������       ��:���D@7             U@
                           @�U�	y�@�           ��@                           �?l�v�]@�           H�@������������������������       ��W��@�             s@������������������������       �,�&�VW@G           p@                           �? {4d�;@�           ��@������������������������       �0���G @�            �l@������������������������       ���+��?@D           �~@                          �<@K��4�@M           ��@                          �7@���{@           ��@                            @� �[l�@d            �@������������������������       �K�=�4@           �y@������������������������       �)��s�@c            �d@                           �?R�����@           �@������������������������       �OƵX�	@           Py@������������������������       �_%Hyg�@           �|@                           �?�~7���@�            u@                            �?:_G�b�@M             _@������������������������       �_j��rd@"            �L@������������������������       �Id�Lҁ@+            �P@                          @A@̫�|�@�            �j@������������������������       ��$�*iD@v            �h@������������������������       ����A�@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     0s@     H�@     �@@      F@     �{@     �U@     ��@     �j@     �@     0y@      =@      @     @^@      r@      *@      1@      j@     �@@     `�@     @U@     �}@     �g@      "@      �?      5@      R@      �?      @      D@             �n@      3@     �b@     �E@      �?      �?      ,@      @@      �?      �?      <@             �Q@      2@     �K@      =@                      @      $@                      $@              C@      @      8@      @              �?      $@      6@      �?      �?      2@              @@      *@      ?@      7@                      @      D@               @      (@              f@      �?     @W@      ,@      �?              @      ;@                      @             �a@             @R@      @                              *@               @      @              A@      �?      4@       @      �?      @      Y@      k@      (@      ,@      e@     �@@     P{@     �P@     �t@      b@       @      @     �P@     �Y@      "@      (@     @]@      9@     `c@      K@      c@      Z@      @       @      :@      D@       @      �?     �G@      .@     �P@      2@     �C@     �H@      �?      @     �D@     �O@      @      &@     �Q@      $@     @V@      B@     @\@     �K@      @             �@@     @\@      @       @      J@       @     �q@      (@      f@     �D@       @              *@      ;@                      $@      �?     �^@      @     �G@      @                      4@     �U@      @       @      E@      @      d@      "@      `@     �A@       @      .@     @g@     �p@      4@      ;@     `m@     �J@     Pr@      `@     pt@     �j@      4@      &@      c@     �k@      .@      0@      g@     �B@     Pp@      Z@     `q@     `b@      4@      @      S@     �[@      @       @     �R@      (@      \@      <@     �S@     @Q@      @      @      M@     �Q@      @       @     �J@      "@      W@      8@     �J@      B@       @              2@      D@                      5@      @      4@      @      :@     �@@      �?      @     @S@     �[@      $@       @     �[@      9@     �b@      S@     �h@     �S@      1@      @      G@      M@      "@      @     �Q@      1@     �D@     �E@      O@     �@@      1@       @      ?@     �J@      �?      @      D@       @      [@     �@@      a@     �F@              @     �@@      F@      @      &@     �I@      0@      @@      8@     �H@      Q@              @      @      :@       @      @      (@      @      ,@      @      4@      9@                      @      0@                       @      @      $@      @      @      *@              @      �?      $@       @      @      $@       @      @      @      .@      (@              �?      ;@      2@      @      @     �C@      &@      2@      2@      =@     �E@              �?      6@      *@      �?      @     �C@      &@      2@      1@      <@      D@                      @      @       @                                      �?      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJnq�6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @I7Q6CA@�	           ��@       	                    �?JLy���@t           6�@                          �5@�Ӑ@	@            D�@                          �2@��Ui�@�           ��@������������������������       ��`�0yv@�            �t@������������������������       �n�B�ض@           py@                          �:@�]<��	@/           ��@������������������������       ����	@U           ��@������������������������       �a�?n�	@�            0u@
                           �?ўj>)8@t           P�@                          �9@�&N�>R@r             g@������������������������       ��GM-�@`            `c@������������������������       ���i<�@             >@                            @����@           y@������������������������       �����.@�            `p@������������������������       ���ʲ��@W            `a@                          �4@�����@9           ��@                           @-�ԍ� @8           ��@                            �?�6�2@�            @j@������������������������       ��߶�p� @,            @S@������������������������       ��Ǹ]��@X            �`@                           �?n�J�̉@�           P�@������������������������       �.XG�H��?�            0q@������������������������       ��K���@
           py@                          �7@�9W]F@           ��@                            �?�D���@�            �x@������������������������       �[�/F�4@�            �j@������������������������       �~_���@r            �f@                           �?lIZ��N@           Pz@������������������������       ���@o            `e@������������������������       �CZ�|`
@�            @o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      r@     ��@      @@     �G@      |@     @V@     `�@     �j@     ��@     �u@      =@      3@      i@     `u@      9@     �C@     �r@     �Q@      w@     �e@     0x@      o@      :@      3@      c@      p@      7@      <@     `n@      K@     @l@     @_@     �p@     �h@      9@       @      M@     @[@      @       @     �W@      (@      c@     �F@     �b@     �T@      @      @      7@      H@               @     �I@       @      T@      1@     �P@     �@@       @      @     �A@     �N@      @      @      F@      $@     @R@      <@     �T@      I@      @      &@     �W@     `b@      0@      4@     �b@      E@     @R@      T@     �]@     �\@      2@      @     @R@     @X@      @      .@     @Z@      3@     �F@      F@     �T@      D@      *@      @      6@      I@      $@      @     �E@      7@      <@      B@      B@     �R@      @             �G@     �U@       @      &@     �L@      1@      b@      I@     �]@      J@      �?              .@      1@                      ,@      @     �N@      &@     �I@      *@                      ,@      .@                      $@      @     �M@      @     �C@      &@                      �?       @                      @               @      @      (@       @                      @@     @Q@       @      &@     �E@      ,@     �T@     �C@      Q@     �C@      �?              8@      @@              $@     �@@      $@     �H@      :@      J@      9@      �?               @     �B@       @      �?      $@      @      A@      *@      0@      ,@              �?     �V@      m@      @       @     �b@      2@     Ѓ@      C@     �z@     @Y@      @              C@     �[@      @      @      F@      @     �x@      3@      k@      J@                      (@     �D@                      @      @      S@      @     �H@      1@                      @      ,@                                      C@      @      $@       @                      "@      ;@                      @      @      C@      @     �C@      "@                      :@     �Q@      @      @     �C@      �?     0t@      (@     �d@     �A@                      $@      8@                      $@             `d@      @      L@      @                      0@      G@      @      @      =@      �?      d@      @     �[@      =@              �?      J@     �^@       @      @      Z@      ,@     `m@      3@     �j@     �H@      @              3@      R@                      G@      (@     �`@      @     �V@      3@      @              $@     �J@                      6@      @     �R@      @      D@      @                      "@      3@                      8@      @      M@              I@      .@      @      �?     �@@      I@       @      @      M@       @     �Y@      .@     �^@      >@              �?      (@      :@                      4@      �?     �B@      $@      J@      (@                      5@      8@       @      @      C@      �?     �P@      @     �Q@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��qhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @E��zC@�	           ��@       	                    �?��-i	@O           ��@                           �?��a-q@�           ��@                           �?�%Mu@�            �r@������������������������       �:��+�@2            @U@������������������������       �t�>]�@�             k@                           �?�nf�S@�            �t@������������������������       ��q�]UH@�             o@������������������������       ����'��@5            @T@
                          �:@u�	���	@�           �@                           �?!Oc~|?	@	           T�@������������������������       ��/��&�	@#           ��@������������������������       ��sie�k@�            0v@                           @O�>�	@�             s@������������������������       ��I���	@.            �Q@������������������������       �9��j�@�            �m@                          �4@
���W@6           ,�@                           @ALP]>X@L           �@                           �?`�?j�=@�             o@������������������������       �8��OKM�?3             W@������������������������       ���,m�@[            �c@                          �0@~j.�4� @�           P�@������������������������       �?���A�?7             U@������������������������       �ɑk+Ϥ @�           ��@                           @���k<@�           @�@                            @�P-{6@<           P�@������������������������       �F��@           �{@������������������������       ��|0q @4            �S@                          �7@~��H@�            �o@������������������������       �`]]053@S            @\@������������������������       �W��/�@[            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �s@     ��@      8@      I@      |@     �U@     ��@      j@     p�@     �v@      <@      6@     @m@     �t@      3@     �C@     �r@     �R@     `v@      f@      u@     @p@      9@             �O@     @W@      @      @     @P@      @      e@      <@      `@     �P@      @              =@      F@      @      @      ;@       @      X@      .@      H@      @@                      @      @                      "@             �B@              6@      @                      6@     �D@      @      @      2@       @     �M@      .@      :@      9@                      A@     �H@               @      C@      @      R@      *@      T@     �A@      @              <@     �C@               @     �B@             �F@      (@     �L@      ;@       @              @      $@                      �?      @      ;@      �?      7@       @       @      6@     `e@     �m@      0@      @@      m@     �Q@     �g@     �b@      j@      h@      5@      "@      `@      j@      $@      >@     �f@      I@     �e@      ]@     �f@     @`@      1@      "@      Z@     �b@      @      8@     `b@     �C@      X@      U@     �[@     @X@      1@              9@      N@      @      @      B@      &@      S@      @@     @R@     �@@              *@      E@      ?@      @       @      I@      4@      2@      @@      9@     �O@      @      @      "@      @      �?      �?      @      @      �?      @       @      2@      @      @     �@@      ;@      @      �?     �F@      ,@      1@      9@      1@     �F@                     �S@     �l@      @      &@     �b@      (@     ��@     �@@     �{@     �Z@      @              A@     �`@      �?      @     �E@      @     �z@      *@     `o@      H@                      2@     �L@                      @      @     �Y@      @     �F@      (@                       @      2@                                      G@              8@       @                      0@     �C@                      @      @      L@      @      5@      $@                      0@     �S@      �?      @      B@             �t@       @     �i@      B@                              5@                                      @@              ;@      @                      0@     �L@      �?      @      B@             �r@       @     `f@      @@                     �F@     �W@      @      @     �Z@      "@     @m@      4@     `h@      M@      @             �A@     �N@              @     @R@      @     �e@      @     �_@      C@      �?              ?@      N@              @     �N@      @     �`@      @     �Z@      B@                      @      �?                      (@      �?      C@              4@       @      �?              $@      A@      @      @      A@      @     �N@      ,@     @Q@      4@       @              @      8@       @              .@       @      >@      �?      9@      "@       @              @      $@       @      @      3@      �?      ?@      *@      F@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJnWhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?ZO�R1@�	           ��@       	                    �?냺w�~@�           t�@                           �?��3���@2           �}@                            @�xۨ��@{            �h@������������������������       �U1�T�@\             b@������������������������       �<��U�X @            �I@                           �?��h}��@�            �q@������������������������       ����I,@Z            @b@������������������������       ��ݧլk@]            �`@
                          �3@U�r��@�            �@                           @/aK( @�            `v@������������������������       �����I@(             Q@������������������������       ��a����?�             r@                          �:@����H!@�            �u@������������������������       ��xY�s�@�            �q@������������������������       ���/�)�@'            �N@                          �4@�q*�@�           X�@                           @|��q @�           ��@                           �?Oj �@�            �h@������������������������       �w�����@/            @P@������������������������       �^O�Ǜ�@V            �`@                           �?�A���@e           ؎@������������������������       �O�
�.A@�            �s@������������������������       ��eƴ"z@�           �@                           @�ߙ� 	@�           (�@                           �?7 |��	@i           Ў@������������������������       �'k�UZ@�             o@������������������������       �鷕��
@�           �@                           �?��p�@c           ��@������������������������       �U�dJ��@�            �q@������������������������       ��-T�z�@�             q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     Ps@      �@      C@      L@     0}@     �U@     $�@      i@     x�@     @v@      9@      �?     �U@     @b@       @      @     �Y@      @     {@      A@     �p@     �T@      @      �?     �H@     @Q@      @      @      O@      �?      Y@      7@     @[@     �H@      @      �?      1@      8@                      6@             �J@      @      L@      0@      @      �?      ,@      1@                      3@             �@@      @     �C@      0@      @              @      @                      @              4@      �?      1@                              @@     �F@      @      @      D@      �?     �G@      3@     �J@     �@@      �?              .@      6@      @      @      4@      �?      :@      ,@      7@      1@                      1@      7@               @      4@              5@      @      >@      0@      �?             �B@     @S@      @       @     �D@      @     �t@      &@      d@      A@      �?              7@      >@              �?      (@             �f@      @     �V@      .@                       @      @                      �?              0@       @      ;@      "@                      .@      9@              �?      &@             �d@      @      P@      @                      ,@     �G@      @      �?      =@      @      c@      @     @Q@      3@      �?              *@      ?@      @      �?      <@      @      `@      @      M@      .@                      �?      0@                      �?              8@      @      &@      @      �?      &@     �k@      w@      >@     �H@     �v@      T@     ��@     �d@     �@     q@      4@      @     �Q@     @d@       @      ,@     �_@      1@      v@      M@     �p@     @Z@      @       @      8@      1@      �?      @      :@       @      I@      *@     �D@      4@              �?      @      @      �?      �?      @              (@      @      6@      "@              �?      5@      &@               @      3@       @      C@      $@      3@      &@              �?      G@      b@      @      &@     @Y@      .@      s@     �F@     �k@     @U@      @      �?      >@     �@@      �?      @      N@      &@     �K@      4@     �I@     �D@      @              0@      \@      @      @     �D@      @      o@      9@     �e@      F@               @      c@      j@      6@     �A@     �m@     �O@     �n@      [@     �q@      e@      0@       @     @]@     �a@      0@      ?@     �c@     �I@     �Y@     �V@     @^@      a@      ,@              1@      D@      �?      (@      H@      @      @@      7@      <@      D@      @       @      Y@     �Y@      .@      3@     @[@     �G@     �Q@     �P@     @W@      X@      &@              B@     �P@      @      @      T@      (@     �a@      2@      d@      @@       @              <@      A@      @      @      I@      @     �Q@      @     @Q@      2@       @               @      @@      @              >@       @      R@      .@      W@      ,@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�^jJhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@Vt0�B@�	           ��@       	                    @�t��qz@�           Ԝ@                          �1@�A[�s@A           @�@                           �?��t�>@�             p@������������������������       �u���=�@k            @e@������������������������       ��G^F]�@4             V@                           �?^,6�X�@�           0�@������������������������       �2^j(RV@           P|@������������������������       � ��n�@�             h@
                            �?�pР�f@V           h�@                           @���H�?�            �l@������������������������       �)Op�� @,             R@������������������������       ��O)#���?f            �c@                          �1@�3���@�           @�@������������������������       �i�d5Jp@�            0q@������������������������       ���Bѻ�@           P{@                          �<@�X��e@<           (�@                           �?x+��@]           $�@                           @�T�[n	@�           x�@������������������������       ��;�(�@o           ؁@������������������������       �a�S�<	@�            �j@                           !@ç(��=@k           Ѝ@������������������������       ����@c           X�@������������������������       ��}W�J�?             .@                            @���%�@�            �t@                           @_N��@�            �j@������������������������       ���C?8h@D            �Z@������������������������       ���fk@K            �Z@                           @�n�#L|@P            �]@������������������������       ���ýK\@C            @Y@������������������������       �;6�|.� @             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     pr@      �@      @@     �P@     |@     �Q@     ��@     �i@     ��@     Pw@      :@      @     @\@     0p@      @      7@     @f@      .@     �@     @U@     �x@     `c@       @      @     �Q@     �a@       @      .@      `@      ,@     �h@     @Q@      e@     �V@      @              4@     �D@                      <@             �R@      4@      F@      >@                      ,@      >@                      9@              ?@      &@     �A@      8@                      @      &@                      @              F@      "@      "@      @              @      I@      Y@       @      .@     @Y@      ,@     @^@     �H@     @_@     �N@      @      @      C@     �Q@              *@     �Q@      (@      S@     �A@     @U@     �F@      @              (@      =@       @       @      ?@       @     �F@      ,@      D@      0@                     �E@     �]@      @       @     �H@      �?     �y@      0@     �k@      P@      @               @      ;@              @       @             �_@      @      E@      1@                      �?      ,@                                      ?@      @      (@      &@                      �?      *@              @       @              X@              >@      @                     �D@     �V@      @      @     �D@      �?     �q@      *@     �f@     �G@      @              $@      C@              @      .@              _@       @     �Q@       @      @              ?@     �J@      @      �?      :@      �?     @d@      &@     �[@     �C@              *@     �f@     �s@      ;@     �E@     �p@     �K@     `w@     �^@     �z@     @k@      2@      &@      c@     �p@      5@     �A@     @l@      G@     pu@     �W@     �w@     @b@      .@      $@     @V@     �_@      1@      7@     �_@      4@     @Y@     �P@     ``@      P@      $@      "@     �R@     @T@      (@      .@     @Y@      0@     �R@      ?@     �[@      E@      @      �?      .@     �F@      @       @      9@      @      ;@     �A@      4@      6@      @      �?      P@     �a@      @      (@      Y@      :@     @n@      =@     �n@     �T@      @      �?      M@     �a@      @      (@      Y@      4@     @n@      <@     �n@     �T@      @              @       @                              @              �?                               @      =@     �H@      @       @     �F@      "@      ?@      ;@      I@      R@      @              7@      :@              @      ;@      "@      .@      ,@     �C@     �J@      @              @      (@              @      ,@       @      $@      @      1@      B@      @              2@      ,@                      *@      @      @      &@      6@      1@               @      @      7@      @      @      2@              0@      *@      &@      3@               @      @      7@      @      @      ,@              $@      *@      @      1@                      �?                              @              @              @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�[2hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?vi�@�	           ��@       	                    �?��+C�@           t�@                           �?r����@�           ��@                            �?���4'�@�             n@������������������������       ��4��@)            @P@������������������������       �����@j            �e@                            �?�ޞ� @           �z@������������������������       ��s9���?A             ]@������������������������       ��u���c@�            �s@
                          �5@�8��ܓ@^           ��@                          �2@�aS [@�            �u@������������������������       ��( �� @k            �e@������������������������       ��&�Ky@h            �e@                           �?e7K�о@�            �l@������������������������       ����X�@N             `@������������������������       �b�.�@=            @Y@                           @ªeb@�           ؤ@                           �?�0ɿ��	@�           �@                           �?���r�	@�           �@������������������������       ��_^�d@            z@������������������������       �hk(�u
@�            �@                           @�Q��@�            �w@������������������������       �6
�a��@2            @S@������������������������       �w蓊F@�            �r@                          �6@1	��O@�           ��@                           �?��x�.@�           H�@������������������������       ���p�L�@            �K@������������������������       ��3��@�           ��@                            �?�E�@�            pv@������������������������       ����n@q             f@������������������������       �K��0=@l            �f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      r@     `�@      >@      I@     `|@     �S@     ��@     �f@     ��@     pt@     �@@             @S@      f@      @      @     �[@      @     p}@      >@     �q@      S@      @              @@     �W@      @      @      O@      @     �p@      1@     `a@     �C@      �?              2@     �C@      @      @      =@      @      L@      (@     �F@      9@      �?              @       @                      (@       @      2@      @      .@      @                      ,@      ?@      @      @      1@      @      C@      "@      >@      6@      �?              ,@      L@               @     �@@      �?     �j@      @     �W@      ,@                              @                      &@              O@              ?@      @                      ,@     �H@               @      6@      �?     �b@      @     �O@      "@                     �F@     @T@                     �H@             `i@      *@     �a@     �B@      @              6@     �H@                      .@             @b@      @     �S@      ;@      �?               @      5@                      &@              W@      @      ;@      "@      �?              ,@      <@                      @              K@       @      J@      2@                      7@      @@                      A@             �L@       @     �O@      $@      @              5@      3@                      :@              7@      @      ;@      @      @               @      *@                       @              A@       @      B@      @              7@     �j@     �y@      9@      F@     pu@     �Q@     p�@     �b@     (�@     `o@      <@      7@     �a@     `p@      3@     �C@      n@      M@     �j@     �_@     �j@     @e@      ;@      7@     �]@     �f@      1@      ?@      h@     �D@     �a@      Y@     �c@     @_@      ;@       @      <@     �Q@      @      &@     �S@      @      P@      ?@      M@      M@      @      5@     �V@     @[@      (@      4@     @\@     �A@     @S@     @Q@     @Y@     �P@      6@              6@     �T@       @       @     �H@      1@      R@      :@     �K@     �F@                      �?      &@              @      .@              ,@      @      @      4@                      5@     �Q@       @      @      A@      1@      M@      4@      I@      9@                     @R@     �b@      @      @     �Y@      *@     �w@      9@     �r@     @T@      �?             �D@      Z@      @      @      K@      "@     �r@      "@     �i@      F@      �?              �?      .@                      @      @      $@              0@      @                      D@     @V@      @      @     �H@      @     0r@      "@     �g@     �C@      �?              @@      G@               @      H@      @      S@      0@     �X@     �B@                      *@      9@               @      $@       @      ?@      &@      O@      5@                      3@      5@                      C@       @     �F@      @      B@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJF�FhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�ѷ]�`@�	           ��@       	                    @c���~@Q           ��@                           �?�,���@�           ��@                          �3@���'�@�            px@������������������������       ��$�X@�            `o@������������������������       �ꀝ��N@J            �a@                            �?2p;��@�           ؄@������������������������       �:�+=L@�             j@������������������������       ���\�@6           �|@
                          �4@�L��J@�           �@                           @`��wѹ@C           X�@������������������������       ��^0W�@!           ��@������������������������       �,k�R��?"             M@                           �?]����@p             f@������������������������       �F�����@)            �Q@������������������������       �Ѹ�Xw&@G            �Z@                            @�v��@I           ��@                           �?���΂�@�           T�@                          �:@�~y���	@J           ��@������������������������       �!��a	@�            �t@������������������������       ����*��@            �h@                           @*+k��-@�           �@������������������������       ���8ƈ�@6           �@������������������������       �t���2@w            �h@                          �=@{Ai(4�@R           ��@                           �?�)m�B@           �{@������������������������       ��P�fR"	@�            �r@������������������������       �qj6���@e            �b@                           �?�a�Td�@8            �U@������������������������       ����sm@             7@������������������������       �����@*             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �s@     @�@     �A@      M@     0}@     �U@     4�@      m@     ��@     �v@      <@      @     @`@     �q@      "@      5@     �k@     �@@     ��@     �U@     �|@      e@       @      @     �S@     @b@      @      2@     �b@      7@     �o@     �P@     �f@     @^@      @             �@@     �A@      �?      �?      F@      �?     @`@      2@      U@      E@       @              2@      3@              �?      8@      �?     �T@      $@      O@      A@                      .@      0@      �?              4@              H@       @      6@       @       @      @     �F@     �[@      @      1@     �Z@      6@      _@     �H@     �X@     �S@      @              ,@      @@                      @@      @     �D@      6@     �@@      ;@      �?      @      ?@     �S@      @      1@     �R@      0@     �T@      ;@     �P@      J@      @              J@      a@      @      @     @Q@      $@      }@      3@     @q@      H@      �?              H@      Z@      @       @     �H@      @     �y@      .@      l@      F@                     �E@      Z@      @       @     �H@      @     Px@      (@      j@     �A@                      @                                              9@      @      0@      "@                      @     �@@              �?      4@      @      J@      @      J@      @      �?               @      4@                      @      @      5@      @      (@                               @      *@              �?      *@      �?      ?@              D@      @      �?       @     �g@     �m@      :@     �B@     �n@     �J@     �s@     @b@     �r@     @h@      4@      @     �]@     `d@       @      <@     @f@      E@     �l@     @Z@     �i@      a@      3@      @      M@     �R@      @      5@     �T@      0@      K@      M@      Q@     �R@      2@       @     �D@      O@       @      .@     �G@      @      ?@     �@@      J@      <@      *@      �?      1@      (@       @      @     �A@      $@      7@      9@      0@     �G@      @             �N@     @V@      @      @      X@      :@      f@     �G@      a@      O@      �?              :@     @R@      @      @      P@      6@     �a@      <@     �X@      G@                     �A@      0@               @      @@      @     �@@      3@      C@      0@      �?      @     �Q@     �R@      2@      "@     @Q@      &@     �U@     �D@      W@     �L@      �?      �?      N@     �O@      *@      @     �J@      &@     �S@      ?@     @V@     �D@      �?      �?     �F@      F@      *@      @     �D@      &@      A@      =@      G@      >@      �?              .@      3@               @      (@             �F@       @     �E@      &@              @      $@      &@      @      @      0@               @      $@      @      0@                              @              �?      @                       @      �?      @              @      $@       @      @      @      $@               @       @       @      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ^�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���n@�	           ��@       	                    �?��[��@!           Г@                           �?)߫�@-           �}@                            @[�@{            `i@������������������������       �{O�Y@Z            @b@������������������������       �������?!            �L@                           �?��#�@�            @q@������������������������       ���eG@S            �`@������������������������       �����@_             b@
                            �?�Q*�@�           ��@                           @�L�ǙZ@v            �g@������������������������       ���j��@9            �V@������������������������       ��,c�N��?=            �X@                           �?���K/�@~           ��@������������������������       ��Y��:�@�            v@������������������������       ��I�L��@�            �n@                           @/��t_@�           ��@                           @�.½X	@�           ��@                           @-��F?(	@V           |�@������������������������       �T)1^u@�           `�@������������������������       �HF��C�	@�           ��@                           �?�zM��G	@            �i@������������������������       �ZBjwi	@[            @c@������������������������       �L�k6�@$            �J@                           @���fg�@�           ��@                           �?��di@           h�@������������������������       ��
�#�@           �x@������������������������       �y�9��@�            �w@                            �?=_ա�@�            �u@������������������������       ��d����@x            �g@������������������������       �����V@]            �c@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     0�@      >@     @Q@      |@     @S@     P�@     �k@     ��@     Pu@     �E@             @T@     `g@      �?      ,@     @\@      1@     �{@      G@     0r@     �P@      @             �B@     �V@      �?      "@     �N@      @     �W@      >@     �Z@     �D@       @              *@      <@                      7@              M@      @     �M@      .@      �?              *@      4@                      5@             �@@      @     �B@      .@      �?                       @                       @              9@              6@                              8@      O@      �?      "@      C@      @     �B@      8@      H@      :@      �?              @      @@      �?      @      5@      @      5@      &@      ,@      (@                      1@      >@               @      1@              0@      *@      A@      ,@      �?              F@     @X@              @      J@      &@     �u@      0@      g@      9@      @               @      6@               @      &@      @     �W@      @      F@      @       @               @      0@               @      @      �?     �C@              8@               @                      @                      @      @     �K@      @      4@      @                      E@     �R@              @     �D@      @     p@      (@     �a@      4@       @              :@     �G@              @      :@      @      c@       @     �S@      "@                      0@      <@                      .@      @      Z@      @      O@      &@       @      2@     �j@     �v@      =@     �K@     �t@      N@     `�@     �e@     ��@     0q@     �B@      1@     `b@      n@      1@     �@@     @m@     �G@     �j@      b@     �l@     �e@      9@      "@     �_@     `i@      0@      ?@      h@     �B@     `h@     �\@     �j@      c@      4@      @     �O@     @X@      @      "@     �[@      8@     �Z@      I@      ^@     @V@      @       @      P@     �Z@      (@      6@     @T@      *@      V@      P@     �W@      P@      1@       @      4@     �B@      �?       @      E@      $@      3@      >@      ,@      3@      @       @      $@      ;@      �?      �?      A@      "@      &@      2@      (@      2@      @              $@      $@              �?       @      �?       @      (@       @      �?              �?      Q@     �^@      (@      6@     @Y@      *@     `u@      >@     �r@     �Y@      (@      �?     �G@     �T@       @      @      N@      @     @q@      1@      j@     @P@      "@      �?      6@      H@              @      C@      @     �a@      @     �V@      C@      "@              9@      A@       @      @      6@      @     �`@      (@     �]@      ;@                      5@     �D@      $@      0@     �D@      @     �P@      *@     �V@      C@      @              *@      6@       @      "@      1@       @      @@       @      L@      ;@                       @      3@       @      @      8@      @      A@      @     �A@      &@      @�t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ|ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��P�@�	           ��@       	                   �;@��~m�E	@�           �@                           �?�f��@D           ��@                           �?5��4X@           `y@������������������������       ��j�/@b            �c@������������������������       ��*���,@�             o@                           �?,�G�4	@B           P�@������������������������       �(�6�*�@�            @w@������������������������       �З� ��	@\           ��@
                           @Z�5��	@�            r@                          �<@�Q�GJj	@�            �o@������������������������       �V�HW�i	@             J@������������������������       �Z�b_%�@|             i@                           �?B��x�@            �B@������������������������       ����c���?             &@������������������������       ���u�}@             :@                           �?�q�;�@�           �@                           �?@20���@�           ��@                          �<@P�����@
           �|@������������������������       �ԜFeZC@           `{@������������������������       �U��2�-@             2@                           @��|��e@�            �t@������������������������       ���_D��?�            �j@������������������������       ���L��@J            @]@                           @b�`��@�           ܗ@                          �5@̨S6�W@�            0x@������������������������       �t�G@@�            @j@������������������������       �g��˻�@p             f@                          �5@]�`���@�           Б@������������������������       �]�LYy@�           H�@������������������������       ��)�6@           �|@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �q@     �@      @@     �J@     �{@     @S@     D�@      i@     H�@     �u@     �@@      0@     @e@      l@      5@      @@     �m@     �H@     �n@      `@     `p@     `g@      :@      $@     �`@     @h@      0@      1@     �i@      ;@     �l@     �X@      n@      ^@      5@             �C@      K@      @      @     �I@      @     @[@      3@     �X@      7@      @              @      0@                      2@             �L@      @      F@       @      �?              @@      C@      @      @     �@@      @      J@      (@      K@      .@       @      $@     �W@     �a@      *@      ,@     @c@      7@      ^@      T@     �a@     @X@      2@              @@     �Q@       @      @     �K@      @      Q@      @@      P@      B@      @      $@      O@     �Q@      &@      "@     �X@      3@      J@      H@     �S@     �N@      ,@      @     �B@      ?@      @      .@     �@@      6@      1@      >@      5@     �P@      @      @      B@      ?@      @      .@      9@      2@      ,@      4@      3@     �O@      �?      @      $@      @       @       @       @      @       @              @       @      �?      �?      :@      :@      @      *@      1@      &@      (@      4@      0@     �K@              �?      �?                               @      @      @      $@       @      @      @                                                       @              @       @       @              �?      �?                               @       @      @      @               @      @      �?     �[@      t@      &@      5@     �i@      <@     ؈@      R@     �@      d@      @              >@      Y@      @       @      G@       @     pv@      ,@     �g@      ?@      �?              1@     @Q@               @      ?@      @      k@      @      V@      4@                      1@     @Q@               @      ?@      @     @j@      @     �U@      1@                                                              @      @       @       @      @                      *@      ?@      @              .@      �?     �a@      "@     �Y@      &@      �?              (@      3@                      "@      �?     @Y@      @      P@      @                      �?      (@      @              @             �D@      @     �C@       @      �?      �?     @T@     �k@       @      3@      d@      4@     @{@      M@     @x@      `@      @              7@      Q@       @      @     �F@      &@     �V@      @@     �Q@      C@      �?              @      D@       @      @      7@      @     �P@      ,@      @@      0@                      1@      <@              �?      6@      @      7@      2@      C@      6@      �?      �?      M@      c@      @      (@      ]@      "@     �u@      :@     �s@     �V@      @              4@      W@      @      @      N@      @     �m@      (@      i@     �D@      @      �?      C@      N@      @      @      L@      @     @[@      ,@     @]@      I@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�1�=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?e��C@�	           ��@       	                     �?I%<�( 	@           ܙ@                           �?��i��@D           �@                           �?	����@f            `c@������������������������       ���B|@-            @Q@������������������������       �;<��@9            �U@                          �:@�!_�Ɗ	@�            �v@������������������������       ��z�u�>	@�            0r@������������������������       ��8�l-@*            @Q@
                          �<@5�j1�@�           Б@                           �? <��]�@z           X�@������������������������       ���z
�@�            `x@������������������������       �"1�Z�
	@�           (�@                            @�g�)s@a             a@������������������������       �^�=(@*            �M@������������������������       ����+	@7            �S@                          �3@����@�           ��@                           @�ov���@J           X�@                           �?|�܋3�@�            `x@������������������������       �Sn���@o             e@������������������������       �ޯc�@�            �k@                           �?�UQw��?X           (�@������������������������       ����8q�?�            pt@������������������������       ��Y��H�?�            �k@                            �?<Ꙛ�@C           ��@                          �5@�t]ˎv@�           �@������������������������       �����@�            @o@������������������������       ��6B�g�@           �|@                           @�mQ�H@�            �@������������������������       ���ڡ�@�            pp@������������������������       ��*�2\@�            �u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Pq@     Ѐ@      8@     �K@     0�@     �U@     �@     �j@     ��@     0w@      >@      2@     �d@     `p@      0@      @@      q@     �K@     �o@     �^@     `m@     �i@      1@      @     �G@     �Q@       @      1@      U@      4@      V@      C@      V@     �I@      @      �?      .@      7@              @      3@       @      B@      @      E@      $@              �?      @      "@              @      $@       @      8@      @      &@       @                      &@      ,@                      "@              (@      �?      ?@       @               @      @@     �G@       @      ,@     @P@      2@      J@      A@      G@     �D@      @      �?      @@      E@       @      *@     �K@      &@      F@      5@      D@      8@      @      �?              @              �?      $@      @       @      *@      @      1@      �?      .@     �]@      h@      ,@      .@     �g@     �A@     �d@     @U@     `b@     @c@      $@      (@      Y@      f@      $@      &@     @e@      @@     @d@     �P@     �`@     �]@      $@      @     �@@     �S@       @      @      L@      @     �R@      :@      L@     �H@              "@     �P@     �X@       @      @     �\@      :@      V@     �D@     @S@     �Q@      $@      @      2@      .@      @      @      2@      @      @      2@      ,@     �A@              �?      "@      @                      @       @      @      @      @      8@               @      "@      &@      @      @      *@      �?       @      *@       @      &@                      \@     @q@       @      7@     �n@      ?@     �@     @V@     `�@     �d@      *@              @@     �X@      �?      @     �N@             �z@      ?@     `n@     �C@      �?              6@     �L@                      6@             �a@      5@     @Z@      5@                      ,@      6@                      (@              J@      ,@      G@       @                       @     �A@                      $@             �V@      @     �M@      *@                      $@     �D@      �?      @     �C@             �q@      $@     @a@      2@      �?              @      :@      �?       @     �@@             �f@      @      P@      $@                      @      .@               @      @             �Z@      @     �R@       @      �?              T@     @f@      @      3@      g@      ?@     Pu@      M@     �q@     �_@      (@             �J@     �V@      �?      @     �U@      1@     @g@      B@     @d@      P@      @              &@      F@              �?      :@      $@     �Q@       @     �Q@      ,@       @              E@      G@      �?      @     �N@      @      ]@      A@      W@      I@       @              ;@      V@      @      (@     �X@      ,@     `c@      6@     �]@     �O@       @              *@     �D@      �?             �H@      *@      L@      .@     �G@      :@       @              ,@     �G@      @      (@     �H@      �?     �X@      @      R@     �B@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJU��HhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @e�)��g@�	           ��@       	                    �?aEg>�@o           ��@                          �;@�c�<	@�           Ę@                           �?�|G�@Q           ̔@������������������������       ������@           �x@������������������������       ��{��=	@M           0�@                            @z�ڵ%�	@�            �o@������������������������       ��9k�g@X             b@������������������������       �W >��@D            @[@
                          �4@�|915@�           `�@                          �3@�l2� U@�             r@������������������������       �62L��@�            `m@������������������������       ��#�t@%            �K@                          �5@��>U@�            �r@������������������������       �m�e;��@"             M@������������������������       �,yX��*@�             n@                          �7@���u%@=           0�@                           @8��O�@@           ��@                          �1@�ְ4�@V           x�@������������������������       �<�O���?�            �q@������������������������       ����4��@�           ��@                          �1@`��Q�i@�            �w@������������������������       ����)@7            �W@������������������������       �����{@�            �q@                           @x��N��@�             z@                           @���_@�            `m@������������������������       �<MS(ѿ@b            �c@������������������������       ��֕��� @0             S@                          �;@�ӊ".N@k            �f@������������������������       ���"�ڞ@G            @_@������������������������       �T���@$             L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�       �@@     �s@     ��@      5@      L@     |@     �R@     �@      m@     x�@     �v@      7@      ?@     �l@     �t@      2@      C@      t@     �J@     Pu@     �f@     pv@     �n@      6@      ?@     �f@     �m@      1@      >@     Pp@      C@     @j@     �`@      m@     `h@      2@      ,@      c@     �i@      *@      8@     �l@      =@     �g@      \@     @j@      a@      .@             �F@     �Q@      @      @     �J@      @     @R@      2@     �U@     �B@       @      ,@     �Z@      a@      "@      3@     �e@      :@     �]@     �W@     �^@     �X@      *@      1@      <@      >@      @      @     �@@      "@      3@      7@      7@     �M@      @      &@      @      "@      �?       @      ;@      @      @      0@      1@      D@      @      @      6@      5@      @      @      @      @      (@      @      @      3@                      H@      X@      �?       @     �N@      .@     ``@      G@     �_@      J@      @              ,@     �I@      �?      @      9@             �T@      9@     �P@      5@                      &@     �C@               @      .@             �Q@      7@      L@      3@                      @      (@      �?      @      $@              (@       @      $@       @                      A@     �F@              @      B@      .@     �H@      5@      N@      ?@      @                      "@              �?      @      @      *@      @      0@      @                      A@      B@               @      ?@      &@      B@      1@      F@      9@      @       @      V@     `p@      @      2@     �_@      6@     h�@      J@     �x@      ^@      �?              O@      j@      @      "@     �S@      *@     h�@      :@     �q@     �S@      �?             �D@     �c@              @      D@      $@     @{@      (@     �h@      G@                      @     �D@                      "@             �c@      �?      N@      @                     �A@     �]@              @      ?@      $@     Pq@      &@      a@      E@                      5@      I@      @      @     �C@      @     @^@      ,@     �V@     �@@      �?              �?      ,@              @      @              :@       @     �@@      @                      4@      B@      @      @     �@@      @     �W@      @     �L@      >@      �?       @      :@     �J@              "@      H@      "@      X@      :@     �Z@     �D@               @      ,@      D@              @      ;@       @     �M@      "@     �O@      0@               @      *@      5@              @      5@       @      A@      "@     �D@      *@                      �?      3@                      @              9@              6@      @                      (@      *@              @      5@      @     �B@      1@     �E@      9@                      @      @              @      (@      @      =@      ,@     �C@      ,@                      @      "@              @      "@      @       @      @      @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJr2!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @��'�Wc@�	           ��@       	                    @y2n?�@�           �@                           �?�)-���@Z           ��@                          �6@y�o)�@           py@������������������������       �z2��:�@�            �o@������������������������       ��q�*��@g            @c@                          �5@=�c8w	@W           �@������������������������       ��/#�ܦ@#           `|@������������������������       ������
@4           �}@
                           �?��g�n@�           ��@                          �6@�2�V@�            �@������������������������       ����Y	 @e           ��@������������������������       �\�sߌ�@~             i@                           @��7]@R@�           ��@������������������������       ��يO_@�           ��@������������������������       ��tc��@             &@                           @@[� g@�           L�@                           �?4�g@��@           ��@                           �?�C$�>	@�            �@������������������������       ��*���R	@|            �g@������������������������       �;�?�	@$            ~@                           �?���@k             f@������������������������       �ɇm�T8@-            �T@������������������������       ��<���@>            �W@                           �?sq�:\r@�            0p@                           @�Ut5b��?8            �U@������������������������       �r[O�l<�?            �A@������������������������       �D�H<�?!            �I@                           @��OvO@o            �e@������������������������       �U��b8@?            �X@������������������������       ��G�w�@0            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@      t@      �@      :@      L@     �|@      S@     �@      m@     �@     �u@      =@      1@     @l@     `w@      *@     �A@     �s@     �J@     ��@     �b@     8�@     �l@      2@      ,@     �a@     �e@       @      ;@     `h@      B@      k@     @^@     �o@      a@      .@              H@     �G@      �?       @      F@      @     �Z@      (@      [@      @@      @              4@      8@      �?      �?      9@      �?     �U@       @     @R@      (@      �?              <@      7@              �?      3@      @      3@      @     �A@      4@       @      ,@      W@     �_@      @      9@     �b@      @@     �[@     @[@      b@     @Z@      (@      @     �B@     �Q@      �?      "@      R@      @     �U@     �E@      U@     �D@      �?      &@     �K@      L@      @      0@     �S@      :@      9@     �P@      N@      P@      &@      @     �U@      i@      @       @     @^@      1@     ��@      >@     �v@      W@      @      @      I@     �Y@       @       @     �T@      @     �q@      *@     �d@      H@       @              =@     �M@       @      @     �P@      @     �o@      @     @Z@      A@      �?      @      5@      F@               @      1@              >@      @     �N@      ,@      �?              B@     @X@      @              C@      (@     p@      1@     �h@      F@      �?              @@     @X@      �?              C@      &@      p@      1@     `h@     �E@      �?              @               @                      �?      �?               @      �?               @     �W@     @e@      *@      5@     �a@      7@     `m@     �T@     @g@     @^@      &@       @      U@     �b@      $@      1@     @_@      6@     �^@     �S@      `@      X@       @       @     @R@     �[@       @      0@     @[@      2@     @T@     �N@      X@      U@       @       @      1@      A@       @      @      9@      @      ?@      (@      8@      ;@      @      @      L@      S@      @      "@      U@      *@      I@     �H@      R@     �L@      @              &@      D@       @      �?      0@      @     �D@      1@      @@      (@                      @      0@       @              "@      @      ,@      @      3@      @                      @      8@              �?      @              ;@      &@      *@      @                      $@      4@      @      @      2@      �?     @\@      @      M@      9@      @               @      @              @       @              K@      �?      2@                                      @                                      :@              @                               @       @              @       @              <@      �?      *@                               @      ,@      @      �?      0@      �?     �M@      @      D@      9@      @              @      @                      &@      �?     �B@      �?      <@      @      @               @       @      @      �?      @              6@       @      (@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ(~�HhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @XIV@s@�	           ��@       	                    �?/;�ڎ�@x           �@                           @�EyL6	@�           �@                           @��O���@�           ��@������������������������       ��O/ZK@�           (�@������������������������       �u�C\�	@�           @�@                            �?��2���	@T            �b@������������������������       ��5�@             J@������������������������       �9�#
�@8            �X@
                           �?���6[@y            �@                          �=@���&�q@w            �f@������������������������       ��}K�}�@p            �d@������������������������       ��KF��P�?             .@                          �3@<����@            y@������������������������       ���{j�@j             e@������������������������       �`TLdm	@�            �l@                           �?Le�%�^@D           �@                           �?�@.��@i           @�@                          �9@�� ��&@�            �s@������������������������       ��9ޱ� @�            �q@������������������������       ��hqaG��?             =@                            �?��Ԝ�L@�            �m@������������������������       �s(!�} @)            �O@������������������������       ��-��C<@s            �e@                            �?߽zV+@�           h�@                           @_���@�           �@������������������������       ��C�X|2@#           p}@������������������������       ���(�g[@}            `i@                          �1@l��qF@;           �@������������������������       ��j���?0            �R@������������������������       �����@           �z@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      s@     ��@      D@      J@     �~@     �S@     ȍ@     �m@     ȉ@     �u@      >@      0@     `i@     �s@      >@     �B@     �t@      M@     `v@      h@     @w@     `n@      <@      0@     �c@     @m@      <@      9@      p@      E@      k@     �a@     p@     @i@      9@      *@      b@     `k@      ;@      8@     �l@     �@@     �i@     @]@     �n@      g@      (@       @     �M@     �Y@      &@       @      X@      *@      Y@      J@     `b@     �S@      "@      @     @U@     @]@      0@      6@     �`@      4@      Z@     @P@     �X@     �Z@      @      @      ,@      .@      �?      �?      <@      "@      (@      9@      &@      2@      *@              "@      @      �?              $@      @              @      $@      @      @      @      @      &@              �?      2@      @      (@      2@      �?      .@      "@             �F@     �T@       @      (@     �Q@      0@     �a@      I@     �\@     �D@      @              1@      .@               @      7@       @      P@      @     �D@      $@                      .@      .@               @      1@       @      O@      �?     �D@      $@                       @                              @               @      @                                      <@      Q@       @      $@      H@      ,@     �S@      F@     �R@      ?@      @              @      <@              @      3@             �K@      5@      >@      "@                      8@      D@       @      @      =@      ,@      7@      7@      F@      6@      @             �Y@     �k@      $@      .@      d@      5@     ��@      F@     P|@      Z@       @              7@      S@              �?     �B@      $@      o@      *@     @`@      *@                      ,@     �D@              �?      8@      @     �c@      @     �N@      "@                      ,@     �A@              �?      8@             `b@      @      J@      "@                              @                              @      $@              "@                              "@     �A@                      *@      @      W@      $@     @Q@      @                              @                      @      @      A@      @      $@      �?                      "@      =@                      @      @      M@      @     �M@      @                      T@     `b@      $@      ,@     �^@      &@     �u@      ?@     0t@     �V@       @             �I@     �R@      @      @      O@       @     @h@      4@     �h@     �L@                      ?@     �J@       @              A@      @      d@      @     �a@      D@                      4@      5@       @      @      <@      @      A@      ,@      L@      1@                      =@     @R@      @       @     �N@      @      c@      &@     @_@      A@       @                      0@                       @              9@              ?@                              =@     �L@      @       @     �M@      @     �_@      &@     �W@      A@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJΎ9KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @%S��O@�	           ��@       	                    �?����@�           n�@                           �?���'O@�           �@                          �<@<f2���@?            @������������������������       ���[��`@           �{@������������������������       �p���@&             M@                           �?�!�܈@o            `e@������������������������       �6x��w@7            �U@������������������������       ��C��d�@8             U@
                          �4@H͌�h�	@�           h�@                           @)5ᦋ=@o           h�@������������������������       �3Z��@e           ȁ@������������������������       ������ @
             4@                          �6@�o_S��	@i           h�@������������������������       ��z�JW1	@�            0q@������������������������       ��wl:��	@�           Ѕ@                          �6@�'�P�@"           H�@                           @5�T��S@�           ��@                            �?)]��	F@�            Pq@������������������������       �fj3�E@,             Q@������������������������       �1��Q�a@�             j@                          �3@�ڰ�R@6           x�@������������������������       �0/q�� @g           @�@������������������������       �f�Ґ�@�            pt@                          �<@6����@@           �~@                           @,��w@           �y@������������������������       ��	&H	�@�            �n@������������������������       ���
�@l            �d@                           �?�����@<            �T@������������������������       ����L@             5@������������������������       �c��^F@-            �N@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     P�@      7@     �I@     �}@     �V@     X�@     `j@     ؈@     @v@      D@      .@     �i@     0t@      5@      D@     pu@     @R@     �w@     �f@     �v@      o@      A@      �?      O@     @R@      �?      @      V@      @     @e@      D@     `c@     @P@      @      �?     �H@     �P@      �?      @      S@       @     @Z@      ?@     �Z@     �J@      @      �?     �E@     �L@      �?       @     �P@       @     �Y@      ;@      Y@      B@      @              @      "@              @      $@              @      @      @      1@                      *@      @               @      (@      �?     @P@      "@     �H@      (@      �?              @      @               @       @      �?      A@      @      2@       @                      @      @                      @              ?@      @      ?@      @      �?      ,@     �a@     @o@      4@     �@@     �o@     �Q@      j@     �a@     �j@     �f@      >@      @     �B@     @W@       @      @     �X@      0@     �\@      L@     �V@      O@      (@      @      B@      W@       @      @     �V@      0@     @\@      L@     �U@      O@      @              �?      �?                      @              �?              @              @      "@     �Z@     �c@      2@      =@     �c@      K@     �W@     �U@     �^@     @^@      2@      @     �B@      F@       @      (@      E@      0@     �E@      8@      ?@      5@              @     @Q@     @\@      0@      1@     �\@      C@      J@     �O@     �V@      Y@      2@             @W@     �l@       @      &@     �`@      2@     ��@      <@     �z@      [@      @              H@     �c@              @      S@      $@     `@      0@     0s@      O@      @              <@      L@                      1@      @     @W@       @      K@      2@      @              @      4@                      �?              2@      �?      1@      @                      8@      B@                      0@      @     �R@      �?     �B@      &@      @              4@      Y@              @     �M@      @     �y@      ,@     �o@      F@      @               @     �J@              @      B@             �q@      "@     �d@      5@       @              (@     �G@              �?      7@      @     @_@      @     �U@      7@      �?             �F@     �R@       @      @     �L@       @     �^@      (@     @^@      G@                     �A@      N@      �?      @      B@       @     �[@      &@     �[@     �A@                      7@      C@              �?      1@      @      T@       @     �O@      3@                      (@      6@      �?      @      3@      @      ?@      "@     �G@      0@                      $@      .@      �?      �?      5@              &@      �?      &@      &@                              @                      @              @      �?      @       @                      $@      $@      �?      �?      2@              @              @      "@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJS��jhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @
�6@�	           ��@       	                    �?|����@d           2�@                           �?Y�0 1	@�           ��@                          �4@n�,�@/           P~@������������������������       �L����!@{             i@������������������������       ������@�            �q@                           @L%���	@�           `�@������������������������       �u�]�ؙ	@o           ��@������������������������       �<P7\=	@R             `@
                           �?	l�m/@t           ��@                          �1@]#��}�@m            �c@������������������������       ���?U1�?            �A@������������������������       ��?�?�@[             _@                           �?��D�9�@           �{@������������������������       ��nOØP@             D@������������������������       ��Q�'S~@�            Py@                           �?�g����@2           ��@                          �5@�9+Of� @k           ��@                            �?Qe6���?           �y@������������������������       �V.�'��?�            @l@������������������������       ���*C��?v            �g@                            @���|x@c            �b@������������������������       �N�C��@T            �_@������������������������       ��<}��?             5@                           �?�I���@�           ��@                           @���h@^           Ё@������������������������       �74��Q@           �z@������������������������       �!�[�%@[            @b@                           @��U̾@i            �@������������������������       ���z��@H             _@������������������������       �|����|@!           �|@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     x�@      B@      N@     �|@     �S@     $�@     `j@     ��@     �u@      =@      1@     `h@     Pt@      8@     �H@     �t@     �N@     �v@      f@     y@     �l@      9@      1@     �c@     �l@      3@      C@     Pp@     �G@      l@     @^@     �q@      f@      9@       @     �H@     �S@      �?      @      Q@             �V@      ;@     @\@     �F@      @               @      :@              @      <@              M@      (@     �I@      &@      @       @     �D@     �J@      �?      @      D@              @@      .@      O@      A@       @      .@      [@     �b@      2@      @@      h@     �G@     �`@     �W@     �d@     �`@      4@      $@     @X@      `@      2@      ?@     @e@      E@     �^@      R@      d@     �]@      (@      @      &@      6@              �?      7@      @      (@      6@      @      *@       @              C@     �W@      @      &@     @R@      ,@     �a@     �K@     @^@     �I@                       @      ,@                      0@      �?      K@      @     �I@      &@                       @       @                                      0@              .@                              @      (@                      0@      �?      C@      @      B@      &@                      >@     @T@      @      &@     �L@      *@     �U@     �I@     �Q@      D@                       @       @               @       @              @      @       @      @                      <@     @R@      @      @     �K@      *@     �T@      F@      Q@     �@@              �?     �U@     @i@      (@      &@      `@      2@     ؄@     �A@     �z@     �]@      @              2@     �Q@      �?      @      4@      @     �q@       @      _@      ;@       @              ,@      I@              @      (@              m@      @     �R@      5@       @              @      >@              �?       @              ^@      @      E@      3@                      &@      4@              @      @             @\@      �?      @@       @       @              @      4@      �?               @      @      J@      @      I@      @                      @      4@      �?              @      @     �B@      @      G@      @                                                      �?              .@      �?      @                      �?      Q@     �`@      &@      @      [@      .@     �w@      ;@      s@     �V@       @      �?     �A@     @Q@      @      @     �L@      "@      h@      ,@     �_@     �J@       @      �?      :@     �G@              �?      F@      @     �c@       @     @V@     �D@       @              "@      6@      @      @      *@      @      A@      @     �B@      (@                     �@@     �O@      @             �I@      @     �g@      *@     �f@      C@                       @      4@      �?              1@      @      =@      @      8@      .@                      9@     �E@      @              A@      �?      d@       @     �c@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��8yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?_��@|	           ��@       	                    �?9�!�&�@s           0�@                           �?�\�pO@           �|@                           �?[�È��@^            �b@������������������������       �R%�l@(            �O@������������������������       ���XS@6            �U@                           �?��Af	@�             s@������������������������       ��6r�"q@K             ]@������������������������       �ܽ���i	@u            �g@
                           �?w �nH$@U            �@                           �?��@�            �p@������������������������       ��'T��?:            @X@������������������������       ��o��`�@h            @e@                           @����@�            �s@������������������������       ��_'
�@@            @\@������������������������       ���;�� @s             i@                          �4@z8��%@	           z�@                          �1@"��L�d@R           4�@                           �?���jY_@           |@������������������������       �XV�U @t            �f@������������������������       ��2�ݘ@�            �p@                           @M�D� @5           `�@������������������������       �#rM��@           @|@������������������������       �C�C@$           �|@                           �?A�GWo0@�           ��@                           �?�}؉�@	           @|@������������������������       �� ډ��@�            @j@������������������������       ��C��@�            @n@                          �9@;�%�O�@�           ��@������������������������       �z��[@�           ��@������������������������       ��V!	@�            �w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �q@     ��@     �@@     �O@     @z@      T@     �@      i@     @�@     Pv@      :@       @      U@      a@      @      &@     �\@      0@     �s@      K@     �g@     �V@      *@       @     �H@     �R@       @      @      Q@      @     �Q@     �C@     @T@      H@      &@              *@      >@                      2@              C@      @      A@      &@      �?               @      $@                      @              0@      �?      .@      @      �?              @      4@                      (@              6@      @      3@      @               @      B@      F@       @      @      I@      @     �@@      A@     �G@     �B@      $@              @      8@                      ,@      �?      5@      $@      ;@      "@      @       @      =@      4@       @      @      B@      @      (@      8@      4@      <@      @             �A@     �O@      @      @     �G@      &@      o@      .@      [@      E@       @              4@      <@               @      E@       @     �W@       @      K@      5@      �?                      @               @      @       @     �N@              0@      @                      4@      9@                     �A@              A@       @      C@      .@      �?              .@     �A@      @      @      @      "@      c@      *@      K@      5@      �?              @      .@              @              @     �D@       @      6@      (@      �?              "@      4@      @              @      @      \@      @      @@      "@              &@     `i@     �z@      ;@      J@     s@      P@     �@     `b@     X�@     �p@      *@      @      J@     �g@      *@      7@     �\@      1@     �}@     �O@     Pr@     �[@      @      �?      5@      O@      �?      @     �A@             `g@      1@     �W@      9@       @               @      2@                      3@              Y@      �?      ?@      @       @      �?      *@      F@      �?      @      0@             �U@      0@      P@      5@              @      ?@     �_@      (@      4@      T@      1@     �q@      G@     �h@     �U@      �?      @      2@      Q@      @      *@      H@      *@     �V@     �A@     @X@     �M@      �?              *@     �M@      @      @      @@      @     �h@      &@     @Y@      ;@              @     �b@      n@      ,@      =@     �g@     �G@     �r@      U@     `r@     �c@      $@              F@     �S@       @      @     �E@      @     �]@      1@     @[@      ?@                      8@     �C@       @      @      3@      �?     �L@      "@     �F@      $@                      4@      D@              �?      8@       @      O@       @      P@      5@              @     �Z@     @d@      (@      8@     `b@      F@     @f@     �P@      g@     @_@      $@      @      M@     �\@      @      0@     �W@      ;@     �a@      <@     @`@     �O@      "@      @     �H@     �G@      @       @     �J@      1@      C@     �C@     �K@      O@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ӭYhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?=>c�-&@�	           ��@       	                    �?�,�Ju�@           h�@                           �?Q��T&�@D           �@                          �:@S��QB@�            �n@������������������������       �(��i�@�            @j@������������������������       ��E�Q�@             B@                          �<@��%��@�            �p@������������������������       ��� ��@�             n@������������������������       �o����Z@             8@
                          �;@�0��$i	@�           p�@                           �?2��H	@H           X�@������������������������       �F�Ճ�	@�            �r@������������������������       ��p�c�@�           ��@                           @���Y�@�             j@������������������������       �d�"9�@M             _@������������������������       �R]�瑊@=            @U@                          �3@aYD���@�           ޡ@                           �?��C�@\           �@                          �0@�����?�             u@������������������������       �7��s��?$            �I@������������������������       �tׁ���?�            �q@                           �?��ҭB@|           h�@������������������������       ���N}M�@�            �p@������������������������       ��L�՘U@�            0t@                           �?n��2h@\           H�@                           @�B�#s@�           0�@������������������������       ��Sn�u@�            q@������������������������       �|Wo'�P@�            Pw@                          �7@�]�}�#@�           `�@������������������������       ����;
�@�            `y@������������������������       �"Su��@�            `s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     @�@      2@      K@     P|@     �S@     �@     �k@     ��@     �v@      :@      3@     `e@     �o@      ,@      >@     �l@      C@      l@     �a@     pq@      j@      2@             �L@     @U@      �?       @      N@      @     @[@      ?@     �[@      E@       @              7@      C@      �?      @      >@      @      M@      7@      C@      ;@                      6@      <@      �?       @      ;@       @      M@      6@      @@      0@                      �?      $@              �?      @      @              �?      @      &@                      A@     �G@              @      >@             �I@       @      R@      .@       @              >@      G@               @      :@             �H@       @     �P@      $@       @              @      �?              @      @               @              @      @              3@     �\@     �d@      *@      6@     @e@     �@@      ]@     �[@      e@     �d@      0@       @     �W@     �`@      *@      4@     @b@      8@     �X@     �V@     @b@      ^@      ,@       @     �A@      O@      "@      @      C@      @      A@      @@      <@      F@       @      @     �M@     �Q@      @      1@      [@      3@     @P@     �M@     �]@      S@      @      &@      4@     �A@               @      8@      "@      1@      4@      7@      G@       @       @      &@      ?@                      "@      @      "@      @      (@      >@       @      @      "@      @               @      .@      @       @      *@      &@      0@               @      `@     �r@      @      8@     �k@     �D@     0�@     �S@      �@     �c@       @             �B@     �Z@       @      @      M@      @     �y@      :@     �l@     �E@      �?              ,@      5@              �?      *@             �f@      @     �V@      &@      �?                       @                      @              <@              @      @                      ,@      *@              �?       @              c@      @      U@      @      �?              7@     @U@       @      @     �F@      @      m@      5@     �a@      @@                      3@      B@      �?              ?@             @Y@      "@      K@      .@                      @     �H@      �?      @      ,@      @     �`@      (@     �U@      1@               @      W@     @h@       @      3@     �d@      C@     �x@     �J@     �q@      ]@      @       @     �E@     �W@      �?      &@     �R@      ,@     �h@      2@     �]@     @P@      @       @      3@      C@      �?       @     �B@      &@     �L@      &@      K@      =@      @              8@     �L@              @      C@      @     �a@      @      P@      B@      �?             �H@     �X@      �?       @     �V@      8@     �h@     �A@     `d@     �I@                      :@      K@               @     �G@      @     �a@      @      X@      9@                      7@     �F@      �?      @     �E@      1@     �J@      =@     �P@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJR�$hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�J��KB@�	           ��@       	                    �?fw����@!           ��@                          �<@j^H��@�           8�@                            �?�,k��@�           �@������������������������       ��ֶU @[            `a@������������������������       �Q�;�O@%           �}@                            �?�s%?@             B@������������������������       �V $UI+�?             &@������������������������       ������@             9@
                           �?����@�           (�@                           �?ӑr�@�            pp@������������������������       ��b�nR@?             W@������������������������       ��mU�В@j            `e@                          �8@���7ay@�            �u@������������������������       ���A+�`@�            �q@������������������������       ���泭�@&            �P@                           @;	�:�'@�           ��@                          �1@ڜ�O#b	@�           D�@                           �?#&�@`            �b@������������������������       ����\�@6            @T@������������������������       ����AD@*            �Q@                           �?�s��=�	@U           �@������������������������       ����M��	@�           ��@������������������������       �)Uil��@�            �t@                          �7@Pm�J��@�           0�@                           �?��t=�@           ؊@������������������������       �z5!�/�@           Pz@������������������������       ����dǀ@           `{@                            �?����4@�            s@������������������������       �qn�.FC@d            `c@������������������������       ���'@_            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     `s@     (�@      6@      E@     �|@     @S@     H�@     @k@     ��@     v@     �B@      �?     @R@     `h@      @       @     �Y@      &@     �|@      H@      q@     �R@      "@      �?     �D@      U@      @      @     �K@      @     �p@      ;@     @]@     �B@      �?      �?      D@     �R@      @      @      K@      @     �p@      :@     �[@      <@      �?      �?      �?      .@              �?      &@       @     �S@      @      7@      @                     �C@     �M@      @      @     �E@      �?     �g@      7@     �U@      8@      �?              �?      $@               @      �?              @      �?      @      "@                      �?      @                                                      @       @                              @               @      �?              @      �?      @      @                      @@     �[@              �?      H@       @     �g@      5@     �c@      C@       @              8@      P@              �?      =@             �H@      &@      L@      9@      @              "@      6@                      @              3@       @      6@       @      @              .@      E@              �?      7@              >@      "@      A@      1@                       @     �G@                      3@       @     �a@      $@     @Y@      *@      @               @     �C@                      *@              _@       @     �S@      &@      @                       @                      @       @      0@       @      7@       @      �?      7@     �m@      x@      3@      A@     0v@     �P@     �@     @e@      �@     `q@      <@      7@     `d@     �l@      (@      <@     @l@      K@      e@     �a@     �l@     @h@      6@              *@      ;@      �?              $@             �E@       @     �@@      0@                       @      0@      �?              @              ,@       @      6@      *@                      @      &@                      @              =@      @      &@      @              7@     �b@     @i@      &@      <@      k@      K@     @_@     �`@     �h@     @f@      6@      7@      ^@     `b@      "@      5@     �c@     �F@     �V@      Z@     �`@      a@      5@              >@     �K@       @      @     �M@      "@     �A@      <@      O@      E@      �?             �R@     �c@      @      @      `@      (@     Pw@      >@     �q@      U@      @             �I@      `@      @      @     �N@      $@     Ps@      *@     �k@      J@      @              ;@      H@       @      @      E@      @      a@      $@     �\@      ;@      @              8@      T@       @      �?      3@      @     �e@      @     �Z@      9@                      7@      =@      @      �?      Q@       @      P@      1@     @P@      @@      �?              .@      6@              �?      7@      �?      @@      "@     �@@      3@                       @      @      @             �F@      �?      @@       @      @@      *@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJJ!hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?+�*�[@�	           ��@       	                    �?�j:�@�           �@                           �?�MΏ�@$           p}@                           �?�T��@v            �g@������������������������       �d	��B@0             Q@������������������������       �F`��@F            @^@                          �7@�NR��@�            �q@������������������������       ��.C���@l            �f@������������������������       ��N���@B            �X@
                           �?�.Z��@�           h�@                          �7@���q�@	           �z@������������������������       �6�[ƠE @�            �u@������������������������       �0yH�c@4            @U@                            �?�{r[ @�            �s@������������������������       ���m"� @k            �f@������������������������       �8���B�?W            �`@                           @i�謷m@�           
�@                           �?��O���	@�           P�@                           �?�b9���	@�           ��@������������������������       �g܋p��@            �x@������������������������       �b�w	
@�           (�@                          �2@�#Df�+@�            @z@������������������������       �C���[@D            @]@������������������������       �Ό��z@�            �r@                           @��Ϋ+@�           đ@                          �1@	����@g           8�@������������������������       ������?c            �c@������������������������       ��5YW�I@           @�@                           �?���i��@X            @a@������������������������       ������~@#            �L@������������������������       �T����k@5            @T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �r@     ��@     �D@      K@     �}@     @T@     4�@     �j@     �@     `v@     �@@             �Q@     �e@      �?      $@     @\@       @     �}@      ?@     �p@      Q@      @             �F@     �Q@      �?      @      R@      @      \@      5@     @W@     �E@      @              2@      7@                      9@             �M@      @      F@      *@       @              @      @                      $@              5@      �?      3@      @                      &@      0@                      .@              C@      @      9@      $@       @              ;@     �G@      �?      @     �G@      @     �J@      0@     �H@      >@       @              3@      =@              �?      7@       @     �G@      @     �B@      4@      �?               @      2@      �?      @      8@      �?      @      (@      (@      $@      �?              :@     �Y@              @     �D@      @     �v@      $@     `e@      9@       @              4@     �K@              @     �@@      @     �k@      @     @S@      .@                      $@     �H@              @      :@      @     �g@      @     �I@      $@                      $@      @                      @              >@      �?      :@      @                      @     �G@                       @       @     �a@      @     �W@      $@       @              @      @@                      @      �?     �Q@      �?     �N@      @       @              @      .@                       @      �?     @R@      @     �@@      @              0@     �l@     �v@      D@      F@     �v@     @R@     ��@     �f@     �@      r@      ;@      0@     �c@     �k@      >@     �@@     �o@     �N@     �h@     �b@      k@     �h@      7@      0@      `@     �c@      :@      :@     �g@     �E@      `@      Z@      c@     �a@      7@       @      :@     �L@      @      (@      P@      @     �R@     �D@      K@     �G@      @      ,@     �Y@     @Y@      5@      ,@      _@     �B@     �J@     �O@     �X@      X@      1@              <@      P@      @      @      P@      2@     �Q@     �F@      P@     �K@                      @      1@                      (@       @     �C@      0@      ,@      &@                      6@     �G@      @      @      J@      0@      @@      =@      I@      F@                      R@     �a@      $@      &@     �[@      (@     �v@      A@      r@      W@      @             �L@     �_@      @      $@     �X@       @     0t@      9@     �p@     @S@      �?              @      *@                      ,@             �T@             �D@      @                      K@     �\@      @      $@      U@       @      n@      9@     @l@      R@      �?              .@      *@      @      �?      (@      @     �C@      "@      7@      .@      @              &@       @              �?      @       @      6@      @      @      @       @              @      &@      @              @       @      1@      @      3@      (@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�]�ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�m7��G@�	           ��@       	                     �?�η;@�           $�@                           �?h��l@2           @@                           @ �ڽ���?i            �d@������������������������       �Ӽ*җ@;             W@������������������������       � ��û��?.             R@                           �?C����@�             u@������������������������       ����kY@N             _@������������������������       ����+�@{            �j@
                           �?)p|@W           T�@                          �2@��^�@           �{@������������������������       ��=��q_@�             m@������������������������       ���a�@             j@                           @@��@K           ��@������������������������       �M���@�            �u@������������������������       ��NW�^@o            �@                           �?�:��b�@            �@                           �?�E�pV�@y           Ђ@                           �?�ˬ��n@�            pq@������������������������       �z�W���@P            �`@������������������������       ��X4�;�@_            @b@                            �?Ȝ��@�            0t@������������������������       �-G���@-            �Q@������������������������       �F�1'��@�            �o@                           @ͬ(�09	@�           ��@                           @��ֻ!	@            ��@������������������������       �v,�&X�	@�            �@������������������������       �rO+��o@&           |@                           !@e�5/0	@�            �h@������������������������       ��!H���@|             g@������������������������       �^�z|�X�?             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `r@     8�@      >@     �O@     �{@     �U@     h�@      i@     ؈@     @w@      8@      @     �V@     �p@      "@      2@     @d@      2@     h�@     @P@     �y@     @d@      @              3@      P@               @      E@      @     @i@      2@     @\@      A@       @              @      9@              �?      @             @T@      �?     �C@       @                      @      ,@              �?      @             �B@      �?      8@      @                              &@                      �?              F@              .@      �?                      0@     �C@              �?      B@      @     @^@      1@     �R@      :@       @              @      1@              �?      3@      @      D@      "@      5@      &@                      *@      6@                      1@      �?     @T@       @     �J@      .@       @      @     �Q@      i@      "@      0@      ^@      ,@     0|@     �G@     �r@      `@      @      @      @@      Q@      @       @     �P@      @     �V@      :@      R@      N@      @      @      1@     �B@      �?      @     �B@             �N@       @      B@      <@              @      .@      ?@       @      @      >@      @      >@      2@      B@      @@      @             �C@     �`@      @       @     �J@      $@     �v@      5@      l@      Q@      �?              3@      M@      @              :@       @     @\@      *@      S@      ;@                      4@     �R@       @       @      ;@       @     �n@       @     �b@     �D@      �?      &@     �i@     �s@      5@     �F@     �q@      Q@      v@     �`@     x@     @j@      2@             �K@     �W@       @      @     @P@      $@     �a@      7@     �a@      M@      @              F@      D@      �?      @     �D@      �?     �@@      ,@      M@     �B@      @              4@      (@      �?      @      2@      �?      .@      &@      ;@      5@                      8@      <@                      7@              2@      @      ?@      0@      @              &@     �K@      �?              8@      "@     @[@      "@     �T@      5@      �?                      (@      �?              $@      @      3@      �?      *@      @      �?              &@     �E@                      ,@      @     �V@       @     �Q@      ,@              &@     �b@     �k@      3@      C@      k@      M@     @j@      \@     �n@      c@      ,@      $@     @`@     `g@      .@      B@      g@     �H@     �g@     @S@     `l@     �`@      "@      "@     �Y@     @`@      &@      >@     �`@     �C@     �R@      O@     �[@     �V@      @      �?      <@     �L@      @      @     �I@      $@     �\@      .@     @]@      F@       @      �?      3@      B@      @       @      ?@      "@      5@     �A@      1@      1@      @      �?      1@      A@      @       @      >@      @      5@     �A@      1@      1@      @               @       @                      �?      @                                      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�J�9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@���^a?@�	           ��@       	                    �?�e	�&f@�           ��@                           �?}HĲ��@^           h�@                           @��|'S@�            �q@������������������������       ����c�@a            �b@������������������������       �a�?b���?S            �`@                           @��o�<@�             q@������������������������       ��v5�@]            �b@������������������������       �he�-���?M            @_@
                          �1@
j�K2�@3           ��@                           @!g�y@�            �v@������������������������       �\m�^�_@m            �e@������������������������       ����`0 @w            �g@                           @�hR�mH@O           X�@������������������������       �j��3�@�            q@������������������������       ��Nu���@�            @o@                           @�D9�b@           L�@                           �?gR���a	@�           ��@                           �?Y�8��=@�            �x@������������������������       �=�}@�$@�            0s@������������������������       �+��@?            �U@                            @�y���	@�           ԑ@������������������������       �GR��A�	@�           �@������������������������       �|+��3�	@           �}@                           �?�g�
�}@J           @�@                            @At~xP@�            �n@������������������������       ��L���@�            �k@������������������������       �D�M3��?             9@                           @��^�?�@�           ��@������������������������       �9���@�            �@������������������������       ���H �@             1@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@      �@      =@      K@     @}@     �S@     ��@     �n@      �@     pu@      7@      @      R@     �g@       @      "@     ``@       @     Ȁ@      R@     �s@      X@      @              8@     �J@              @      D@             0p@      *@      `@      B@      �?              &@      <@               @      4@             �a@      @     �K@      1@                      "@      2@                      .@              L@      @      @@      .@                       @      $@               @      @             �U@      �?      7@       @                      *@      9@              �?      4@              ]@      @     @R@      3@      �?              &@      (@              �?      .@             �F@       @      G@      1@                       @      *@                      @             �Q@      @      ;@       @      �?      @      H@      a@       @      @     �V@       @     `q@     �M@     �g@      N@      @      �?      ,@     �Q@      �?      �?      <@      �?     �_@      0@     �R@      >@              �?      $@     �D@      �?      �?      0@      �?      D@      0@      9@      4@                      @      =@                      (@             �U@             �H@      $@               @      A@     �P@      �?      @     �O@      @     �b@     �E@      ]@      >@      @       @      4@      ;@      �?      @     �F@      @     @R@      C@      A@      3@      @              ,@      D@              �?      2@      �?     �S@      @     �T@      &@              2@     �j@      v@      ;@     �F@     u@     �Q@     �}@     �e@     `~@     �n@      2@      0@     �d@     �j@      5@     �B@      n@     �K@     �i@     �a@      o@     @f@      0@              H@      F@      @       @     �J@      @     @W@      >@      S@     �@@      �?             �F@     �B@      @      @      G@             �I@      8@     @P@      >@      �?              @      @              @      @      @      E@      @      &@      @              0@      ]@      e@      2@      =@     `g@     �I@     �[@     �[@     �e@      b@      .@      @     @R@      V@      @      5@      Y@      B@     @Q@     �O@      \@     @V@      @      "@     �E@     @T@      (@       @     �U@      .@      E@      H@     �N@      L@      $@       @     �I@     �a@      @       @     @X@      .@     0q@     �@@     �m@     @Q@       @               @      J@       @              8@      @     @X@      @     �D@      .@                       @      J@       @              7@      @     @S@      @      C@      ,@                                                      �?              4@              @      �?               @     �E@     @V@      @       @     @R@      &@     @f@      =@     �h@      K@       @       @      E@      V@      @       @      Q@      @      f@      ;@     `h@      K@       @              �?      �?                      @      @       @       @      �?                �t�bub�     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �1@�)Y�<@�	           ��@       	                    �?��|}�?@y            �@                           �?t�IC�@h            �b@                          �0@��5�?\@.             P@������������������������       �`_`C@             4@������������������������       �mfz1�@!             F@                           @���Y�@:            �U@������������������������       ��%�G��@             E@������������������������       �q  �}l@            �F@
                           �?�N����?           �z@                            @To�r	��?s            �e@������������������������       ��\�m��?Z             a@������������������������       �����?            �C@                           @�g�@�            �o@������������������������       �)�o���?            �A@������������������������       ����@�            `k@                          �8@r�}�#�@           
�@                           �?&V�TN�@�           �@                           @_�DL��@E           ��@������������������������       ��~�h@_           0�@������������������������       �ܸ�{	@�            �v@                           �?�*0:(E@�           ��@������������������������       �a� �z@"           `{@������������������������       �ϫx8=8@d           �@                           @D�A�q	@Q           ��@                            @΋�0��	@�           ��@������������������������       ��U2�!	@�            �w@������������������������       ����w�	@�             l@                            �?`��Y[�@�            `s@������������������������       �����g�@m             e@������������������������       �&Ё}��@[            �a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �p@     Ȃ@     �A@     �N@     �{@     @T@     @�@      m@     @�@     `u@      5@       @      *@      U@       @      @      A@             @o@      5@     �a@      =@               @      @      ;@       @      �?      5@              B@      @     �@@      1@                      �?      @                       @              6@      @      .@       @                      �?                              @              "@      �?       @      @                              @                      @              *@       @      *@      @               @      @      4@       @      �?      *@              ,@       @      2@      "@                      @      .@                      @              &@      �?      @      �?               @      �?      @       @      �?      "@              @      �?      *@       @                      @     �L@              @      *@             �j@      0@      [@      (@                      �?      1@              �?      @              [@             �C@      @                              *@              �?      @             @V@              ;@      @                      �?      @                      �?              3@              (@       @                      @      D@               @      "@             �Z@      0@     @Q@      @                       @      �?                      �?              0@      "@      @                              @     �C@               @       @             �V@      @     �O@      @              *@      p@     (�@     �@@     �L@     �y@     @T@     p�@     `j@     ؅@     �s@      5@       @      g@     �w@      3@     �B@     s@      H@     x�@     @\@     x�@     �g@      &@      @      Z@      d@      "@      8@     `d@      3@     �_@     @P@     @e@     �V@       @      @     �O@     @Z@      @       @     �X@      &@     @V@      7@     �_@     �G@       @      @     �D@     �K@      @      0@      P@       @      C@      E@      F@      F@      @      �?     @T@     �k@      $@      *@     �a@      =@      }@      H@     Pv@     �X@      @              8@     @P@      �?      @      5@      @     �g@      @     �Z@      .@              �?     �L@     �c@      "@      $@     @^@      8@     q@      E@     @o@     �T@      @      @     @R@     �`@      ,@      4@     �Z@     �@@     �_@     �X@     �e@      _@      $@      @      N@     �X@      (@      $@      R@      ?@      Q@     �S@      R@     @V@      $@       @      >@     �M@      @      �?      I@      :@     �D@     �I@      H@      O@      "@      @      >@      D@       @      "@      6@      @      ;@      <@      8@      ;@      �?              *@     �A@       @      $@     �A@       @     �M@      3@      Y@     �A@                      &@      ;@              �?      *@       @      >@      *@      I@      6@                       @       @       @      "@      6@              =@      @      I@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��\thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @����Y@�	           ��@       	                     �?�xB,��@{           ��@                           �?��iQ�V@�           ؃@                           �?q�O��@|            �h@������������������������       ��0g@5             T@������������������������       ���W�@G            �]@                           �?/���j�@           @{@������������������������       ��dH���@N            �_@������������������������       ��yin��@�            `s@
                           �?R�A���@�           @�@                          �<@r�Y:��@'            }@������������������������       ��_ːN@           z@������������������������       �Gqa	_@!            �H@                           @��v.&o	@�           ��@������������������������       ����	(	@s           ��@������������������������       ���R^1	@T             a@                           �?0h۱<�@;           ��@                          �>@Q3>`� @h           �@                            �?<I�Lmt @_           ��@������������������������       ��1ݵ�)�?G            �Z@������������������������       �V	�P1� @           `z@������������������������       �j{��0J@	             *@                            �?�����@�           ��@                          �5@�v�{s@�            �o@������������������������       �t�u�%�@a            �b@������������������������       ���rc/�@J            �Z@                          �<@O�?#>@(           �@������������������������       ���L���@           x�@������������������������       ��/C��n@             �I@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     �s@     ��@     �D@     �M@     �{@     �Q@     ȏ@      k@     P�@     �v@      <@      0@     �m@     `u@      >@     �D@     �r@     �M@     �w@     �f@     �x@     `n@      9@      @      S@      Y@       @      @     �T@      4@     �]@     �J@     �[@      J@      $@      @      ;@      =@                      4@      �?      L@      @     �H@      "@       @      @      @      &@                      "@      �?     �A@      �?      *@      @                      7@      2@                      &@              5@       @      B@      @       @      �?     �H@     �Q@       @      @      O@      3@     �O@      I@      O@     �E@       @              @      1@              @      9@      @      9@      $@      =@      @       @      �?     �E@      K@       @      @     �B@      ,@      C@      D@     �@@     �C@      @      (@     `d@     @n@      <@     �A@     �k@     �C@     Pp@      `@     �q@     �g@      .@             �K@     �K@      �?      $@     �J@      @     �]@      ?@     �W@     �E@      �?             �H@      J@      �?      @     �F@      @     �\@      9@     @V@      =@      �?              @      @              @       @              @      @      @      ,@              (@      [@     `g@      ;@      9@      e@     �A@     �a@     @X@     @g@     �b@      ,@      @     @X@     �d@      ;@      7@      b@      @@     �_@     �Q@     �e@     @a@      &@       @      &@      4@               @      7@      @      1@      ;@      (@      $@      @             �S@     @k@      &@      2@     `a@      &@     �@      B@      x@      _@      @              0@     �R@       @      @      5@      @     �q@      &@     �Z@      6@      �?              0@     �R@       @      @      2@      �?     pq@      "@     @Z@      3@      �?                      ,@       @               @      �?      O@              1@       @                      0@      N@              @      0@              k@      "@      V@      &@      �?                      �?                      @       @      �?       @      �?      @                     �O@     �a@      "@      ,@     �]@       @     Pv@      9@     �q@     �Y@       @              0@      >@                      6@       @      Y@       @     �L@      4@                      @      4@                      *@             �Q@      @      <@      "@                      *@      $@                      "@       @      >@      @      =@      &@                     �G@     @\@      "@      ,@      X@      @     p@      1@     �k@     �T@       @             �A@     @[@      "@      *@     @S@      @      p@      0@     �k@     �Q@       @              (@      @              �?      3@              �?      �?       @      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ԑchG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @��>�XL@�	           ��@       	                   �<@���~��@`           B�@                          �2@��4=�@�           ��@                           �?b�}�@3           P~@������������������������       ��+��|v@�            �u@������������������������       ��6b@^            @a@                           �?���mh5	@�           �@������������������������       ���5��	@�            �@������������������������       ��nN#@�            Px@
                           �?<ԅ�:@�            �n@                          �=@�<�r@1            �V@������������������������       ������.�?             G@������������������������       ��،J@            �F@                          �=@ޑ5۠@b            �c@������������������������       �����,@             G@������������������������       ��;{��@F            �[@                           @bxe @A           ��@                           �?ZB��K�@�           ̒@                          �2@�$6�A @           �{@������������������������       ��5,{�?}            @h@������������������������       ��S�;�	@�            `o@                          �4@%��~��@�           ��@������������������������       ���TX��@�            �x@������������������������       �y���@�            �v@                           @���f@B           P@                            �?�Dݯ@4           �}@������������������������       ��6�ވG@A            @Y@������������������������       �z�R@�            Pw@������������������������       ��~@             ;@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        2@     �p@     x�@      ;@     �J@     �z@      T@     t�@     �m@     Ї@      x@      D@      1@     �h@     �s@      0@      G@     �r@     @P@     y@     �g@     �v@     0q@      <@      *@     `e@     �q@      0@      D@     �p@     �J@      x@     �c@     Pu@     �i@      :@              ?@     @P@              @      O@      @     �a@      >@     �U@     �L@      @              8@     �D@              @     �J@      @     @X@      6@      K@      G@      @              @      8@                      "@      �?      G@       @      @@      &@              *@     �a@     �k@      0@     �B@     �i@      H@      n@      `@     �o@     �b@      7@      *@     �[@     �c@      0@      <@     �c@      B@     @c@     �X@      f@      ]@      7@              =@     �O@              "@      H@      (@     �U@      =@     �S@      A@              @      9@      ?@              @      ?@      (@      1@      ?@      4@      Q@       @               @      @              @      &@               @      $@      *@      >@       @              @       @                      @                      �?      $@      :@                      @      @              @       @               @      "@      @      @       @      @      1@      9@              @      4@      (@      "@      5@      @      C@              �?      @       @              �?       @      @       @      &@      �?      1@              @      *@      7@               @      2@      @      @      $@      @      5@              �?     �R@     @n@      &@      @     @`@      .@     `�@     �H@     y@     @[@      (@      �?      D@     @e@       @      �?     �V@       @     �@      <@     �q@     �P@      @      �?      *@      P@              �?      4@      @     �m@      @     @U@      $@                      @      6@                      @             �a@      �?      6@                      �?       @      E@              �?      0@      @     �X@      @     �O@      $@                      ;@     �Z@       @             �Q@       @     �p@      5@     �h@      L@      @              &@     �J@                      3@      �?     �d@      $@      [@      ;@                      0@     �J@       @             �I@      �?     �Y@      &@     @V@      =@      @             �A@      R@      "@      @      D@      @      b@      5@     �]@     �E@      @              9@     �Q@      "@      @      D@      @     �a@      1@     �\@      E@      �?              @      $@      �?              @      �?     �E@      �?      ;@      @                      3@     �N@       @      @     �A@      @      Y@      0@      V@     �A@      �?              $@      �?                               @      �?      @      @      �?      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��rhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?���KS@�	           ��@       	                    �?3j*�J@           �@                            @����:�@3            @                          �;@�/t12@�            0r@������������������������       �U� Ql@�            �p@������������������������       ��T�}
@             8@                          �=@���@            �i@������������������������       ���g��U@s            `g@������������������������       ���F�z� @             4@
                          �>@�̕2Қ@�           ��@                          �1@ �	 @�           ��@������������������������       �#�N��"�?k            @d@������������������������       ��W�n��@Z           ��@������������������������       ��=W�p@             :@                          �5@��_�,>@�           �@                          �1@�\t�@r           �@                           �?la�G@�             x@������������������������       �>�1/�i@C            @[@������������������������       ��]9.o�@�            0q@                           @�"��]�@�           ��@������������������������       �p(*�g"	@]           `�@������������������������       �{+�š@$            }@                          �;@��3�0	@)           ,�@                           @c���@X            �@������������������������       ��6���@l           Ё@������������������������       ���YT/3@�            `x@                            @ek�2ݫ	@�            �t@������������������������       ����@�            �j@������������������������       ���Z��	@G            @]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        .@     �r@     �@      :@      K@     �~@      T@     ��@     @k@     x�@     �x@      ?@              R@      e@      �?      $@     �Z@      (@     P{@     �C@     pr@     �Q@      @              G@     �U@      �?      "@     �Q@      @     �Y@      6@     @\@      E@      @              8@      F@      �?      @      D@      �?     �L@      (@     �T@      6@      @              5@      D@      �?       @     �B@              L@      (@      T@      .@      @              @      @              @      @      �?      �?               @      @                      6@      E@              @      ?@       @     �F@      $@      ?@      4@                      5@     �B@               @      6@       @      F@      $@      ?@      2@                      �?      @               @      "@              �?                       @                      :@     �T@              �?      B@      "@     �t@      1@     �f@      =@      @              :@     �S@              �?      @@      @     �t@      &@     �f@      7@      @               @      (@              �?      @             �X@              E@      �?       @              8@     �P@                      =@      @      m@      &@     @a@      6@      �?                      @                      @       @      @      @       @      @              .@     @l@     �w@      9@      F@     �w@      Q@     ��@     `f@     �|@     @t@      9@      @     �T@     �h@      *@      1@      e@      :@     @x@      R@     0q@     @c@      @      �?      3@      K@      �?       @      @@              a@      1@     �V@      ?@              �?      *@      &@      �?              2@              5@      @      5@      2@                      @     �E@               @      ,@              ]@      (@     @Q@      *@              @     �O@     �a@      (@      .@      a@      :@     `o@     �K@      g@     �^@      @      @     �B@     �R@      "@      *@      W@      5@     @Y@      H@     �R@     �R@      @              :@     �P@      @       @      F@      @     �b@      @     �[@      H@      �?      "@      b@     �f@      (@      ;@     �j@      E@     @g@     �Z@     �f@     @e@      2@       @     �X@     �a@      "@      .@     �c@      <@     `c@      U@     �a@     @]@      ,@      �?      M@      Q@      @      (@      V@      7@     �V@     �@@     @Y@     @U@      @      �?      D@      R@      @      @     �Q@      @      P@     �I@     �C@      @@      @      @      G@     �D@      @      (@      L@      ,@      ?@      7@     �D@     �J@      @      @      ?@      8@      �?      @     �E@      "@      0@      (@      <@      C@       @              .@      1@       @      "@      *@      @      .@      &@      *@      .@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJw�UhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����Ba@�	           ��@       	                    �?�r�$$�@f           \�@                           @ U��@           0�@                           �?./K4��@d           �@������������������������       �D�w��@�             v@������������������������       �l�o&��@�            �o@                           �?�OG�uB	@�            Pr@������������������������       �����@2            �T@������������������������       ���dz�}	@�            `j@
                           �?�����@N           ��@                          �;@&����)@�            �v@������������������������       �FZFW'{@�            @t@������������������������       ��H��_@             C@                           �?2g�߅	@h           ��@������������������������       �PRz9��	@�           p�@������������������������       �/eF��@�             n@                          �7@=Y���@0           l�@                           �?���Td�@:           <�@                           �?�Ƿ��& @B           �~@������������������������       ��xdX��?�            `q@������������������������       �rRh���?�             k@                            �?���%�@�            �@������������������������       �Gë�\8@m            �f@������������������������       �r���Y@�           P�@                           @G����Z@�            �x@                            �?��g���@�            �k@������������������������       ���)�r�@E            �[@������������������������       �G~�Ꮕ@H            �[@                            �?��.���@i            �e@������������������������       ��`
��U@:             X@������������������������       �<�ڳ@/            �S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �s@     ��@      9@      K@     @|@     �X@     H�@     `l@     ��@     �u@      6@      7@     �l@     Pu@      3@      C@     �s@      S@     w@      g@     @w@     �m@      4@      @     �Y@      a@      (@      .@     �`@      A@      c@     �S@     �_@     @X@       @      �?      K@      W@      "@      @     �V@      :@     @`@      @@      Y@     �P@      �?              B@     �I@      @      @      F@      @     �X@      5@     �K@      A@      �?      �?      2@     �D@      @             �G@      5@      @@      &@     �F@     �@@               @     �H@     �F@      @      "@      F@       @      7@     �G@      :@      >@      @              ,@      (@              @      5@               @      "@      @      "@               @     �A@     �@@      @      @      7@       @      .@      C@      6@      5@      @      4@     �_@     �i@      @      7@     @f@      E@      k@     @Z@     �n@     �a@      (@              ?@     �P@               @     �@@      �?     @S@      &@     �Y@     �A@       @              9@     �M@              �?      <@      �?     @S@      @     @X@      <@       @              @       @              �?      @                      @      @      @              4@     �W@      a@      @      5@      b@     �D@     `a@     �W@     �a@     �Z@      $@      4@     �R@     �V@      @      1@      ]@     �@@      U@     @R@     @[@      V@      $@              5@     �G@      @      @      =@       @     �K@      5@      A@      2@                     �U@     `k@      @      0@     `a@      6@     ��@     �E@     �y@     �[@       @             �P@     �f@      @      $@     �T@      &@     Ѐ@      2@     @s@     �R@       @              *@     @V@              �?      6@      �?     �n@      $@     �Y@      $@                       @      G@              �?      0@      �?     �a@      �?     �K@      @                      @     �E@                      @             �Y@      "@      H@      @                     �J@     �V@      @      "@     �N@      $@     @r@       @     �i@     @P@       @              0@      ,@               @      4@             @T@      �?      C@      $@                     �B@     @S@      @      @     �D@      $@     `j@      @     �d@     �K@       @              5@     �C@       @      @      L@      &@     �W@      9@     �Z@      B@                      &@      8@              @     �C@      @     @P@      @      L@      $@                      @      4@               @      $@      @      @@      @      9@      @                      @      @              �?      =@             �@@      @      ?@      @                      $@      .@       @      @      1@      @      =@      3@      I@      :@                       @      @              @      @      @      1@      "@      ;@      3@                       @      "@       @              *@      �?      (@      $@      7@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJF,/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@��פm@�	           ��@       	                   �1@}ॐ��@\           �@                           @c7mWQ@�           �@                            �?�gw�d@�            �q@������������������������       ���r�$v@Z            �_@������������������������       ���6� @`            `c@                           @�
�W�@�            @t@������������������������       ��R	,ig@�            `r@������������������������       ����k�h@             >@
                           �?��,ڵ@�           ��@                            �?��F�@g           ��@������������������������       ��CT��M@_            �b@������������������������       ���34	@            z@                          �4@Q���v�@s           ��@������������������������       ��.�,]K@�            �@������������������������       �{k)x0c@�            �i@                            @�č'"�@Q           �@                          �<@)Y�]�@           P�@                           @$0��&@�           ��@������������������������       ��sh$C	@k           ��@������������������������       ��+�æ�@           pz@                            �?q�-�u@�            �n@������������������������       �"��o�@u            `j@������������������������       ��{�,�@            �A@                           �?w�(8��@E           �~@                          �=@�����	@�             s@������������������������       ���|a�	@�             p@������������������������       �.���VT@              G@                           �?�4�[;�@y            �g@������������������������       ������@%             L@������������������������       �XI���/@T            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     x�@      @@      H@     p}@     �T@     �@     �p@     ȉ@     �u@     �A@      @     @^@     �r@      1@      5@      o@      6@     ؄@     �Y@     p@     �d@      *@              8@     @R@      @       @     �J@      �?     �o@      6@     @a@      A@      �?              (@      3@              �?      5@             @a@      $@     @P@      ,@      �?               @      (@              �?      (@              N@      @      ;@      "@                      $@      @                      "@             �S@      @      C@      @      �?              (@      K@      @      �?      @@      �?      ]@      (@     @R@      4@                      "@     �J@      @              ;@             �Y@      &@      R@      1@                      @      �?              �?      @      �?      ,@      �?      �?      @              @     @X@      l@      ,@      3@     �h@      5@     �y@      T@     �v@     @`@      (@      @      J@     �R@      $@      &@      X@      "@     �R@      G@      [@     �Q@       @               @      6@               @      >@      �?      4@      ,@     �@@      0@      @      @      F@     �J@      $@      "@     �P@       @     �K@      @@     �R@      K@      @             �F@     �b@      @       @      Y@      (@      u@      A@     p@      N@      @              E@     @\@      @      @     @Q@      @     �q@      =@     �h@      J@                      @      B@              �?      ?@      @     �J@      @     �N@       @      @      @     �f@     �l@      .@      ;@     �k@     �N@     �r@     �d@      t@      g@      6@      @      ^@     @d@      @      6@      d@     �D@     �i@     �Z@     �o@      a@      0@      @      U@     �`@      @      4@      _@      8@     `g@     �T@     �k@      V@      *@      @      O@      S@      @      1@     @U@      1@     �S@     �L@      Z@     �I@      (@      �?      6@     �M@      �?      @     �C@      @     @[@      9@     �]@     �B@      �?      �?      B@      ;@               @      B@      1@      4@      9@      >@     �H@      @      �?      @@      9@               @      6@      .@      0@      8@      ;@      F@      @              @       @                      ,@       @      @      �?      @      @              �?      N@      Q@      "@      @      O@      4@     @V@     �L@     @Q@      H@      @      �?      F@     �F@       @      @      E@      2@      ?@      E@      =@     �@@      @              B@     �A@      @      @      =@      1@      <@      E@      <@      <@      @      �?       @      $@       @       @      *@      �?      @              �?      @                      0@      7@      �?              4@       @      M@      .@      D@      .@                      @      @                               @      6@      $@      $@      @                      *@      1@      �?              4@              B@      @      >@      (@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��[�u@�	           ��@       	                    �?��߄��@
           �@                           �?Q��RD@,           P~@                            �?j��^1=@�            �k@������������������������       ���?�{@C            �[@������������������������       �ާ��Qo@B             \@                          �;@�-��@�            `p@������������������������       ��ه>3�@�             l@������������������������       ���Z��@             C@
                           �?F�g���@�            �@                           @ف��;T@           �{@������������������������       �F�xR�@q            �g@������������������������       �Q�$� !�?�            p@                          �8@�wT�O@�            r@������������������������       ����Z<@�             o@������������������������       ��Ho&�z@            �D@                          �5@�Β��_@�           �@                            @�i��@q           ��@                           @�5��@�           ��@������������������������       �߲��<@r           �@������������������������       �T�|���@           0{@                          �1@+�!���@�            @w@������������������������       ��Wf���@:             Z@������������������������       �=@,d1*	@�            �p@                            �?����T	@8           h�@                          �6@�^c�	@�             u@������������������������       ����@"            �J@������������������������       ��i�[z�	@�            �q@                           @e��9-	@X           P�@������������������������       ��J���	@n           ��@������������������������       ��mi�e@�            �w@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �q@     x�@      =@      O@     �|@     �W@     ��@     @l@     ؈@     �v@      <@       @      Q@     �e@      @      "@     @]@      *@     �z@      C@     �q@     �S@      @       @     �E@     @T@      @      @      P@      @     �W@      8@     �Z@     �J@      @       @      0@      @@      @      @      >@      @      F@      2@      D@      <@               @      @      3@                      ,@      �?      3@      @      5@      6@                      "@      *@      @      @      0@      @      9@      (@      3@      @                      ;@     �H@               @      A@              I@      @     �P@      9@      @              3@     �F@                      =@              H@      @      N@      .@      @               @      @               @      @               @      �?      @      $@                      9@      W@      �?       @     �J@       @      u@      ,@      f@      :@       @              ,@     �L@               @     �A@      @     @k@      @     @W@      2@                      (@      ;@               @      ,@      @     �R@      @     �E@      $@                       @      >@                      5@       @     �a@      �?      I@       @                      &@     �A@      �?              2@      @     �]@      "@      U@       @       @              &@      ?@      �?              ,@             @\@      @     @P@      @      �?                      @                      @      @      @       @      3@      @      �?      3@      k@      x@      9@     �J@     �u@     �T@     ��@     �g@      �@     �q@      7@      @     �Q@     �i@      $@      8@      b@      <@      w@     �V@     0s@      _@      @       @     �G@     @c@      @      ,@     �W@      3@     `r@      O@     �m@     @U@      @       @      ;@      Z@       @      @     �M@      3@     �^@      M@     �]@     �M@       @              4@      I@      �?      "@      B@             `e@      @     @]@      :@      �?      @      8@     �I@      @      $@     �H@      "@      S@      <@     �Q@     �C@      @              @      *@      @       @      @              @@      $@      8@      @              @      1@      C@      @       @     �E@      "@      F@      2@     �G@     �@@      @      (@      b@     �f@      .@      =@     @i@      K@     �g@     �X@     �i@     �c@      1@       @     �G@     �B@      @      (@     �F@      4@      J@      B@     �D@      B@      @      �?      .@      @       @       @      @      @      *@      @              @              �?      @@      ?@      �?      $@      D@      1@     �C@     �@@     �D@     �@@      @      $@     �X@      b@      (@      1@     �c@      A@     @a@      O@     �d@     �^@      (@      $@     �P@     �Y@      &@      &@     @Y@      >@      G@      F@     @S@     �T@      &@              ?@     �D@      �?      @      L@      @      W@      2@     �U@     �C@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�is-^@�	           ��@       	                    �?�
�!:�@           ,�@                           �?�@x�k�@!           |@                            �?��� @j            �d@������������������������       ��e�c�/@H             [@������������������������       ����@"             L@                           �?�w?�15@�            �q@������������������������       �kl��7�@O            �\@������������������������       �njȿ@h            @e@
                           �?��x@�           P�@                          �3@k��<@           �z@������������������������       �qn�) @�            �j@������������������������       ��T,���@�            `k@                            @l%��C@�            �u@������������������������       ��5�W�o@�            Pr@������������������������       �p.�<�?%             K@                          �5@ڿ�ŗG@�           ��@                          �1@��jM��@�           �@                           @�cB�>@�            �v@������������������������       �E�L���@�            �t@������������������������       �����@             9@                           �?͒��)@�           H�@������������������������       �@���?*	@           @x@������������������������       �x�l��@�           p�@                            �?{	)cp	@           �@                           @XSw��	@�            Pw@������������������������       �-'���	@�            @s@������������������������       �0�W	@%            @P@                           @C��J%	@6           x�@������������������������       �j��gL]
@w            �j@������������������������       ���rsg@�           Ѕ@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     q@     ��@      C@     �D@     �}@     �X@     0�@     `l@     �@     pu@     �B@      @     @P@     �e@      @      @     �]@      &@     P{@      G@     r@     �P@      @      @      =@      T@      @      @     �P@      @     �Y@      ;@     �V@      B@      @      @      $@      6@                      8@              I@      @      A@      (@       @      @       @      ,@                      $@              @@      @      6@      (@       @               @       @                      ,@              2@       @      (@                              3@      M@      @      @      E@      @      J@      4@     �L@      8@      �?              $@      3@      @      @      ,@      @      8@      &@      .@      $@                      "@     �C@                      <@              <@      "@      E@      ,@      �?              B@      W@      �?       @     �J@       @     �t@      3@     �h@      ?@      @              2@     �J@               @     �A@      @     @i@      &@     �U@      0@                       @      7@              �?      "@             @\@      @     �F@       @                      $@      >@              �?      :@      @     @V@      @      E@       @                      2@     �C@      �?              2@      �?     �`@       @     �[@      .@      @              2@     �A@      �?              0@      �?     @\@      @      V@      .@      @                      @                       @              4@      @      7@                      *@      j@     �x@      ?@      B@     0v@     �U@     ��@     �f@     �@     @q@      ?@      @     �O@      k@      @      .@     �e@      >@     Pw@     @R@     0s@     �_@      *@              6@      J@      �?      @      =@      �?      `@      ,@     @T@      <@                      5@      J@      �?      �?      7@             �^@      ,@      S@      9@                      �?                       @      @      �?      @              @      @              @     �D@     �d@      @      (@     @b@      =@     �n@     �M@     @l@     �X@      *@      @      ;@      H@       @      $@     �T@      0@     �K@     �A@      N@     �C@      $@              ,@      ]@      @       @      P@      *@     �g@      8@     �d@     �M@      @      "@      b@     @f@      8@      5@     �f@     �L@     �g@      [@     �i@     �b@      2@      �?     �F@     �F@       @      $@      E@      2@      N@      H@      H@      E@      @      �?     �B@      E@      @      $@     �C@      ,@      K@      C@      D@      =@      �?               @      @      @              @      @      @      $@       @      *@      @       @      Y@     �`@      0@      &@     @a@     �C@      `@      N@     �c@      [@      (@      @      7@      9@      &@      @      =@      *@      .@      6@     �E@      3@      @      @     @S@      [@      @      @     @[@      :@     @\@      C@     �\@     @V@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�f�<hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�y��q@�	           ��@       	                    �?}p'8m	@           ��@                           �?)�xK�@2           �}@                           �?��]Ȓ@z            �f@������������������������       ������F@6            �S@������������������������       �m@v�L|@D            @Z@                            �?����l�@�            `r@������������������������       �v����@9            @X@������������������������       ���3�@            �h@
                           �?�T� �	@�           @�@                           @�����@           �y@������������������������       �&��� @;             W@������������������������       ��,��@�            t@                          �2@���UL
@�           ��@������������������������       ���o"˙@K            �`@������������������������       ��+�8�
@�           x�@                          �3@l�"S�@�           ��@                           @5��bs@K            �@                           @�c��@�           ��@������������������������       ���3�@�             v@������������������������       ��	�� �?�            �w@                           @D%�2�M@z            �h@������������������������       ��?S,�@U             b@������������������������       �&�B�@%             J@                           @9~~y�n@U           �@                          �4@���u�@�            �u@������������������������       ��HՅ+;@'            �M@������������������������       ��'!���@�             r@                           @h�%Zb�@~           �@������������������������       ���R{�@�           ��@������������������������       �6&���@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     0r@      �@     �@@      N@      z@     �X@     ,�@     @n@     ��@      v@     �@@      ,@     �e@      p@      2@      E@     �j@     �K@      o@     `c@     `o@     �g@      <@      �?      G@     �R@      @       @     �H@       @     �]@      =@      Y@     �E@       @      �?      *@      <@                      4@             �M@       @      E@      &@      �?      �?      @      $@                      $@              ;@      @      1@      @                      "@      2@                      $@              @@      @      9@      @      �?             �@@     �G@      @       @      =@       @      N@      5@      M@      @@      �?              "@      5@               @       @              0@      $@      9@      @                      8@      :@      @      @      5@       @      F@      &@     �@@      :@      �?      *@      `@     �f@      .@      A@     �d@     �J@      `@     �_@     �b@     @b@      :@              :@     @S@      �?      .@     �K@      ,@     �P@     �A@     �O@      K@      @              @      $@      �?      �?      ,@      @      "@      *@      8@       @       @              4@     �P@              ,@     �D@      $@      M@      6@     �C@      G@      @      *@     �Y@      Z@      ,@      3@     �[@     �C@      O@     �V@      V@      W@      4@              (@      5@       @              :@      �?      *@      (@      8@      2@      @      *@     �V@     �T@      (@      3@      U@      C@     �H@     �S@      P@     �R@      1@      �?      ]@      t@      .@      2@     �i@     �E@     ��@     �U@     �@     `d@      @              A@      ]@      @      @      M@      @     �x@      @@     �l@      G@                      ;@     @X@       @      �?      <@      @      u@      9@      f@     �A@                      0@     �J@                      0@      @     �`@      5@     @V@      5@                      &@      F@       @      �?      (@             `i@      @     �U@      ,@                      @      3@       @      @      >@             �N@      @     �K@      &@                      @      .@       @              2@             �J@      @     �D@      @                      �?      @              @      (@               @      �?      ,@       @              �?     �T@     �i@      &@      *@     @b@      D@     @x@     �K@     `q@     @]@      @              :@     �K@      @      @     �H@      4@      S@      ?@     �J@      ;@      �?              �?      &@      @       @      ,@      �?      .@       @      @      @                      9@      F@              @     �A@      3@     �N@      =@      I@      4@      �?      �?      L@     �b@       @      @     @X@      4@     �s@      8@      l@     �V@      @      �?      3@      ]@      @      @     �O@      ,@     �n@      3@     `d@     �Q@                     �B@     �@@      @      �?      A@      @     �P@      @      O@      3@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJؗ�-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@�����a@�	           ��@       	                    @�(ad6�@v           ̜@                           �?a�I���@D           Ѝ@                           �?E	k�@�           �@������������������������       �.#'"3@�            @r@������������������������       ��xǾ	@�            �u@                           �?yp`�@�            ps@������������������������       ��Ϋ}c�@E            �\@������������������������       �B+ �@v            �h@
                           @�A"�8@2           ȋ@                           @��w�8@�           �@������������������������       �@���//@�            �g@������������������������       �w@�� @%           0~@                           �?h�����@�             k@������������������������       �;��޻f@9            �V@������������������������       �7F)�[@S            @_@                           @}��˅o@)           ,�@                           �?*sS�U	@:           $�@                           �?���$�@�            �t@������������������������       �A����@�            �o@������������������������       � ~i7�a@1            �T@                          �:@��Z��	@`           ؍@������������������������       �m!x?	@�           @�@������������������������       ��|��O�	@�            0s@                          �7@т��Q
@�           h�@                          �6@�VC��@�            �v@������������������������       �~����@�            Pp@������������������������       �{�oc��@D             Z@                           @3�{�܅@            z@������������������������       �y�ǋ��@p            �d@������������������������       �@ŠI�@�            `o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ;@      r@     ��@      =@      P@     @}@     �R@     @�@     �k@     h�@     w@      8@       @     �Y@      o@      $@      @@     @h@      2@     ��@     �P@     �w@     �b@       @       @      Q@      b@      @      3@     �a@      .@      k@      K@     `e@      [@      @       @     �J@     �V@      @      (@     �Z@      ,@     @a@      @@     �Y@     �S@      @      �?      3@     �E@              @      I@      @     �S@      .@     �J@      9@              @      A@     �G@      @      @      L@      &@      N@      1@     �H@      K@      @              .@      K@      �?      @      A@      �?     �S@      6@     @Q@      =@                      @      8@      �?      �?      3@              6@      @      7@      *@                      &@      >@              @      .@      �?     �L@      .@      G@      0@                      A@      Z@      @      *@      K@      @     �y@      *@     @j@      E@       @              7@      U@      �?      @      =@       @     @t@      $@     `d@      @@                      ,@      D@                      "@       @      T@      @     �A@      @                      "@      F@      �?      @      4@             �n@      @      `@      9@                      &@      4@      @       @      9@      �?      U@      @     �G@      $@       @              @      @              @      @             �E@      @      1@      @       @              @      .@      @       @      4@      �?     �D@              >@      @              3@     @g@      t@      3@      @@      q@     �L@     pw@      c@      y@     `k@      0@      1@     �`@     �g@      .@      <@      g@      F@     �e@      _@     �j@      c@      *@      �?      E@      K@      @      @      B@      �?      O@      7@     @S@      =@      �?      �?      A@      I@      @      @      A@      �?      @@      2@      J@      5@      �?               @      @                       @              >@      @      9@       @              0@      W@      a@      (@      7@     �b@     �E@     �[@     @Y@      a@     �^@      (@      @      L@      \@      @      2@     �Y@      <@     �S@      O@     �Y@     @Q@       @      (@      B@      8@      @      @      G@      .@     �@@     �C@      A@      K@      @       @      J@     @`@      @      @     @V@      *@     @i@      =@     @g@     �P@      @              6@     @R@       @              A@      $@     �\@      @      T@      5@       @              (@     �D@      �?              ?@       @     �T@      @     @P@      .@       @              $@      @@      �?              @       @      @@      @      .@      @               @      >@     �L@       @      @     �K@      @      V@      6@     �Z@      G@      �?       @      �?      =@       @      @      ,@      �?     �B@      &@      G@      2@                      =@      <@                     �D@       @     �I@      &@      N@      <@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @Y�Ėxr@�	           ��@       	                    �?���O�@�           ��@                           �?�
����@W           ��@                           �?�9�\X@�            �s@������������������������       �G�]k�!@[            `c@������������������������       �����o@e            `d@                            �?D���'�@�           ȃ@������������������������       �Sc���@v            �f@������������������������       �܉(h�@!           0|@
                          �4@��zY+�@�           0�@                           @r(k8Z@           Ȉ@������������������������       �����@�             t@������������������������       ���7��@/           �}@                           @_����@�           ��@������������������������       �gxg��@1           (�@������������������������       ��4aNn	@Z            �a@                          �1@�"	��s@�           �@                           �?�3��@^            �d@                          �0@���M#@2            �V@������������������������       ��_X��[@             7@������������������������       �ih���@&            �P@                           �?̪� @,            �R@������������������������       � ˬ��~�?             =@������������������������       ��.rn�?             G@                          �?@W^,�i�@]           �@                           �?�#���@F           ��@������������������������       �#��u�@�             r@������������������������       ��9��hp	@�           ��@                           @1��^@             G@������������������������       ��0%�*@
             4@������������������������       ����K�@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     X�@      @@     �M@     �|@      U@     h�@     �h@     (�@     �w@      A@       @      k@     �v@      2@     �B@     �s@     �K@     �@     @`@     ؂@     �o@      7@       @      P@     �`@      @       @     �U@       @     pt@      8@      k@      S@      @       @      @@     �J@       @      �?      E@      @      L@      ,@     �R@      @@      @       @      (@      :@       @              2@      @      @@      (@      :@      3@       @              4@      ;@              �?      8@              8@       @      H@      *@      @              @@     �T@       @      �?      F@      @     �p@      $@     �a@      F@      �?              @      3@       @              ,@       @     @W@      �?     �A@      *@                      =@     �O@              �?      >@       @     @f@      "@     �Z@      ?@      �?      @      c@     �l@      ,@     �A@     @l@     �G@     �y@     �Z@     0x@      f@      0@              J@     �V@      @       @      X@      @     �o@     �@@     �e@      T@      �?              <@      B@       @       @      M@      @      N@      :@      L@      H@      �?              8@     �K@      @      @      C@              h@      @      ]@      @@              @     @Y@      a@      "@      ;@     @`@      F@     �c@     @R@     �j@      X@      .@       @     @T@     �\@      "@      :@     �\@      =@     �a@     �J@     �h@     �V@      $@      @      4@      6@              �?      0@      .@      2@      4@      0@      @      @      1@     �X@      d@      ,@      6@      b@      =@     �p@     �P@     @i@     @_@      &@              0@      ,@       @      @      &@             �S@       @      3@      *@                      $@      $@       @      @      $@             �B@      @      @      @                      @      @              @       @               @      �?               @                      @      @       @               @             �A@      @      @      @                      @      @                      �?              E@      @      (@      @                      �?      @                      �?              0@              @       @                      @                                              :@      @      @      @              1@     �T@     @b@      (@      3@     �`@      =@     �g@     �M@     �f@      \@      &@      (@     �S@     �a@      "@      3@      ^@      =@     �g@     �M@      f@     �Y@      &@              4@     �G@      �?      @      =@             �S@      ,@     �P@      :@              (@      M@     �W@       @      (@     �V@      =@     �[@     �F@     �[@      S@      &@      @      @      @      @              *@                              @      $@              @       @      @       @              @                              @      @               @      @      �?      �?              $@                               @      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ}��/hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�dN�@�	           ��@       	                    �?�����@           "�@                           �?o|ZB�@F           �@                            �?�ٳ�.�@�            pr@������������������������       ��A�;@]            �c@������������������������       �u�Z��@[             a@                           @�����@�           Ѓ@������������������������       ����� @2           �~@������������������������       �g��?@\            �a@
                           �?���@�           ��@                           @CY-��@            `�@������������������������       �Ǽ��M@�           8�@������������������������       �&2�Q]B@@            @Y@                           @����z@�           �@������������������������       �I�7�L@�           ��@������������������������       ��Ғ>Zl@            �A@                           �?y*u�`@�           ��@                           @D���@�            `s@                           �?qQ�,�<@�            `k@������������������������       ��Uc�?            �G@������������������������       �#RԦ@u            �e@                          �3@aK-ZB=�?A            �V@������������������������       �2xajW�?             F@������������������������       ���I�?#            �G@                           @m�LUh�@�           �@                          �9@6���bS	@           ��@������������������������       �Rm����@*           �|@������������������������       �Y$3zh	@U            �a@                           @�x�2�@k            �d@������������������������       �rKAę@>             Y@������������������������       ��� ��@-            �P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �s@     ��@     �A@     @P@     @|@      N@     |�@     �j@     8�@     `u@      6@      @      k@     �z@      6@     �C@     �r@     �G@     (�@      d@     ȁ@     `l@      (@             �Q@     �a@      @      @      T@      @     �u@      9@     @h@     �J@      @              ?@     �G@       @      @     �F@       @     �M@      0@      N@      <@       @              *@     �A@                      9@       @     �B@      @      ?@      $@                      2@      (@       @      @      4@              6@      $@      =@      2@       @             �C@      X@      �?      �?     �A@       @     0r@      "@     �`@      9@      �?              A@     �O@                      4@      �?     @n@      @     �Y@      8@                      @     �@@      �?      �?      .@      �?     �H@      @      @@      �?      �?      @     @b@      r@      3@     �A@     �k@     �E@     p|@     �`@     pw@     �e@      "@      @     @Q@     ``@      @       @      \@      *@     �e@     �P@     �b@     @R@      @      @     �I@     @^@      @       @      Z@       @     @d@      F@     @a@     @P@      @              2@      $@       @               @      @      *@      6@      *@       @       @      �?     @S@     �c@      *@      ;@     @[@      >@     �q@     @Q@      l@     @Y@      @      �?      Q@     �c@      *@      ;@      Z@      ;@     `q@     �P@     �j@     �X@       @              "@      �?                      @      @       @       @      "@       @       @      $@     �X@     �d@      *@      :@     �b@      *@     @o@     �K@     �e@     �\@      $@              6@      C@              @      =@      �?     �\@      .@      N@      9@                      4@     �@@              @      ;@      �?     �N@      ,@     �A@      8@                               @                                      7@      �?      (@      @                      4@      9@              @      ;@      �?      C@      *@      7@      5@                       @      @               @       @             �J@      �?      9@      �?                       @                              �?              8@              1@                                      @               @      �?              =@      �?       @      �?              $@      S@     �_@      *@      4@     �^@      (@      a@      D@     �\@     �V@      $@      $@     �P@     �[@      *@      2@     �X@      &@     �S@     �B@      S@     �S@       @      @      B@      V@      "@      ,@     @V@       @     @Q@      <@      O@     �I@      @      @      >@      7@      @      @      "@      @      "@      "@      ,@      ;@      @              $@      0@               @      8@      �?      M@      @      C@      (@       @              @      @                      1@      �?     �D@              :@      �?       @              @      $@               @      @              1@      @      (@      &@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ_�"hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?�3�/�]@�	           ��@       	                    �?��M	!6	@�           d�@                           �?��&Y�@1           �}@                            �? ��|j�@�             k@������������������������       �	*��,@@O             ]@������������������������       ��[�\O@?             Y@                           �?�)����@�            pp@������������������������       ��M�;-@=            �X@������������������������       ��$�� @f            �d@
                           @b|�!t�	@�           �@                           �?r�N/�	@�           \�@������������������������       ��˚yc�@           �y@������������������������       �s�N N
@�           Ѕ@������������������������       ��ǣ�Ɖ@            �A@                          �3@�N���@�           �@                           �?���ˡ@d           ��@                           @��`�� @�             w@������������������������       ��\?Q�<�?�            �p@������������������������       ��i�H��@>            �Y@                            �?�d��Rp@p           x�@������������������������       ���0Ж)@\             b@������������������������       ��-i�5�@           �{@                            @��E��g@U           Ĕ@                           !@���rf@�           h�@������������������������       ���T=@�           ,�@������������������������       ���*|���?             .@                           @����R@�            pq@������������������������       �0�`@F            �Y@������������������������       ��-v�a�@k             f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        1@     `s@     P�@      >@      M@     �}@      W@     ��@     �i@     `�@     �u@      :@      1@      f@      o@      5@      F@      p@     �G@     �j@     �\@     q@     `h@      4@             �L@     �Q@      �?       @      O@      @     �U@      2@     �\@     �L@                      6@      6@      �?       @      B@      @     �C@      *@     �E@      <@                      &@      $@      �?      @      3@              5@      $@      5@      3@                      &@      (@              @      1@      @      2@      @      6@      "@                     �A@     �H@                      :@             �G@      @      R@      =@                      "@      3@                      @              9@      �?      ?@       @                      :@      >@                      5@              6@      @     �D@      5@              1@     �]@     @f@      4@      B@     @h@     �E@     �_@      X@     �c@     @a@      4@      ,@     @\@     �e@      4@      B@     `g@      E@     �_@     �V@     `c@      a@      .@              ;@      R@      �?      2@     �R@      @     �Q@      >@     �L@      L@              ,@     �U@     �Y@      3@      2@      \@      B@      L@      N@     �X@     @T@      .@      @      @      @                      @      �?              @      @      �?      @             �`@     s@      "@      ,@     @k@     �F@     �@     @W@     ؁@     �c@      @             �G@      `@              @     �M@       @     `w@      ?@     �p@     �E@      �?              5@      A@              �?      2@             `e@      @     �Y@      .@      �?              *@      9@                       @             `a@      �?     �Q@      $@                       @      "@              �?      $@              @@      @     �@@      @      �?              :@     �W@              @     �D@       @     `i@      ;@     �d@      <@                       @      2@              @      "@              Q@      @      B@      @                      8@     @S@               @      @@       @     �`@      7@      `@      7@                     �U@      f@      "@       @     �c@     �E@     �v@      O@      s@     @\@      @              Q@      c@      @      @     �^@     �C@     `q@     �G@     �n@     �T@      @             �P@     �b@      @      @     @^@      >@     `q@     �G@     �n@     �T@      @              �?      @                       @      "@                                                      3@      7@      @       @      B@      @     @U@      .@      N@      ?@      �?              (@      .@      �?              &@       @      2@      (@      0@      0@                      @       @       @       @      9@       @     �P@      @      F@      .@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�h�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @RhJ��\@�	           ��@       	                   �;@����w�@]           �@                           �?�m�-_@�           p�@                          �3@�-����@�           ��@������������������������       ���ٿ��@�            Pq@������������������������       �ܒ��l,	@            |@                          �5@a�	�@�           �@������������������������       �4E[O@�           ��@������������������������       ����0@�@5           �~@
                           �?��g�
@�            pr@                           @��:�!@K            �Z@������������������������       ��v,�.�@=            �U@������������������������       �.Դ��@             4@                           �?�B݋�
@y            �g@������������������������       ��/j��@            �E@������������������������       ������
@_            @b@                          �4@�`UtgH@D           �@                           �?����N�@I           �@                           @>qMP�@9           �~@������������������������       ���K��	@�            �y@������������������������       �5��}�@:            @T@                           @MoJBP�@           `{@������������������������       �F!�,:� @H            �\@������������������������       ��)�g;J@�            @t@                            @=�:11@�           (�@                          �7@�/0w%N@�            �@������������������������       ��|��<@�            �t@������������������������       ���y7C�@�            `u@                           @�?o��A@Q             `@������������������������       �I��{�@J            �\@������������������������       ���
�Q,@             ,@�t�b��
     h�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@     ��@      =@      M@     @}@     �U@     ��@     @j@     8�@     �w@     �A@      .@      k@     Ps@      4@     �F@      s@     �M@     �w@     �e@     �v@     �p@      ;@      @     �f@     @q@      .@      A@     pp@     �C@     @v@     @b@     �t@      j@      9@      �?     �R@     @Z@      @      2@     �Y@      3@      a@      L@     @Z@      W@       @      �?      5@      B@                     �A@      @     �P@      :@      J@     �@@      �?             �J@     @Q@      @      2@      Q@      *@     �Q@      >@     �J@     �M@      @      @     �Z@     `e@       @      0@      d@      4@     `k@     �V@     �l@      ]@      1@       @     �G@     �T@       @       @      W@       @     �c@     �F@     �b@     �O@      "@      @      N@      V@      @       @      Q@      (@      O@     �F@     �T@     �J@       @      "@     �A@     �@@      @      &@     �E@      4@      8@      <@      ;@      M@       @       @      "@      4@              @      0@       @      @       @      &@      8@              �?      @      4@              @      &@       @      @      @      @      4@              �?       @                              @                      @      @      @              @      :@      *@      @       @      ;@      (@      3@      4@      0@      A@       @              (@       @                      "@              @      "@      @       @      �?      @      ,@      &@      @       @      2@      (@      .@      &@      (@      @@      �?             �U@     �k@      "@      *@     @d@      ;@     �@      B@     �y@     �\@       @              D@      ^@      @      @      I@      @     �z@      ,@     `k@     �E@                      1@     �M@      @      @     �A@             �l@      $@     �[@      8@                      (@      K@      �?       @      =@              h@       @     �X@      (@                      @      @      @      �?      @             �A@       @      (@      (@                      7@     �N@              @      .@      @     �h@      @      [@      3@                       @      7@                       @      @     �J@              5@       @                      .@      C@              @      *@             @b@      @     �U@      1@                     �G@     �Y@      @      @      \@      6@      k@      6@     @h@     �Q@       @              F@      W@      @      @      X@      6@      f@      5@      c@      N@      @              2@      J@       @              I@      *@      Y@      @     �R@      .@      @              :@      D@      �?      @      G@      "@     @S@      0@     �S@     �F@                      @      $@       @       @      0@             �C@      �?     �D@      &@      @              �?       @               @      0@             �B@      �?     �C@      &@                       @       @       @                               @               @              @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�%+#hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �? �4R@�	           ��@       	                    �?�ǵ-K�@           ��@                            �?����E�@5           P~@                          �;@/�K�[@[            �`@������������������������       �Z[�[@M             \@������������������������       ���z��@             5@                           �?h| �@�             v@������������������������       ���妨|@M            �]@������������������������       ����K=L@�             m@
                          �>@����-@�           �@                          �3@T�f�Y�@�           ��@������������������������       �����&��?�            @u@������������������������       �p��Q��@�            �u@������������������������       �/p3O�@             .@                           @�ji;/@�           F�@                           @��Jng	@�           �@                           �?IAS��@�           ��@������������������������       ��r��f	@S            �^@������������������������       �1{E��.@t           ��@                           �?*IS��	@           x�@������������������������       �®��3A
@v            �@������������������������       �����]�@�            �i@                            �?kj�@�           t�@                          �6@@��}��@�           �@������������������������       �w,B:�@           �}@������������������������       �fY[���@|            �h@                          �9@݇(D@@            �@������������������������       ��&�t�1@           0y@������������������������       ���0�M�@>            @[@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@     @r@     �@      A@      J@     �}@     @P@     ؎@     @l@     ��@     �v@      ?@      �?     �T@      c@      @      &@     �[@      @     0z@     �B@     `q@      V@      @      �?     �I@      R@       @      @      P@       @     �[@      7@     �W@     �K@      @      �?      (@      ?@               @      &@      �?      7@      @      A@      (@       @              $@      7@               @       @              7@      @     �@@      @       @      �?       @       @                      @      �?                      �?      @                     �C@     �D@       @      @     �J@      �?      V@      3@     �N@     �E@      �?              (@      0@                      $@             �D@      @      >@      @                      ;@      9@       @      @     �E@      �?     �G@      .@      ?@     �B@      �?              ?@     @T@      �?      @      G@      @     @s@      ,@     �f@     �@@                      <@     @T@      �?      @      D@       @     0s@      &@     �f@     �@@                      .@      8@              @      &@             `d@      @     �Z@      *@                      *@     �L@      �?       @      =@       @      b@      @      S@      4@                      @                              @      �?      �?      @      �?                      3@     @j@     �z@      ?@     �D@     �v@      N@     ��@     �g@     �@     Pq@      <@      3@     �a@     �p@      9@      ?@     �m@     �G@     �h@     `c@     �j@     @g@      6@      "@     �K@     �]@      &@      ,@      `@      6@     �V@      L@     @\@     @Z@      @      @      $@      1@               @      4@      @      @      4@      &@      5@       @      @     �F@     �Y@      &@      @     @[@      2@     @U@      B@     �Y@      U@      �?      $@      V@     @b@      ,@      1@     �[@      9@     �Z@     �X@      Y@     @T@      3@      $@     �P@      Y@      *@      1@      U@      4@     �P@     �R@     �Q@     �P@      3@              5@      G@      �?              :@      @      D@      8@      =@      .@                     �P@      d@      @      $@      `@      *@     0w@      A@     `r@     �V@      @             �C@      X@       @       @      K@      $@     �j@      3@     `f@     �H@      �?              6@     �P@       @      @     �A@      @     `f@      @      ]@     �A@      �?              1@      >@              �?      3@      @     �@@      ,@     �O@      ,@                      <@     @P@      @       @     �R@      @     �c@      .@     �\@      E@      @              4@      O@      �?             �E@      @     `a@      @      W@      @@      @               @      @      @       @      ?@              4@      "@      7@      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJnLLhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @� �L41@�	           ��@       	                    �?(����@j            �@                           �?�q�^�	@�           Ę@                            @�>���@0            }@������������������������       �Zf4�@�             o@������������������������       �讝�@�             k@                          �:@|�ދ	@�           |�@������������������������       ����z$	@*           0�@������������������������       �'I�o�	@�             o@
                           �?Z�02�@s           x�@                          �8@1ZR���@k            �e@������������������������       ���� �@W            �a@������������������������       �G�!�y�@             >@                          �5@�Z7��@           0z@������������������������       ���D���@�            @l@������������������������       ��c�y4@}             h@                          �7@_�~j5@M           $�@                           @Xk.��@W            �@                           @�{ǂ�@�            �q@������������������������       ����T� @�            �f@������������������������       ���c�f�@7             Y@                           @�&�NZ@�           ��@������������������������       �E8h8j4 @�           ��@������������������������       �m\<���@�            Py@                            @���ab@�            �x@                          �<@A��ʐ�@�            `t@������������������������       �e�9L=I@�            �o@������������������������       �/��7ע@)            @R@                           @����d@+            �P@������������������������       �D�����?             A@������������������������       ����wx�@            �@@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �t@     0�@      6@      J@     ~@      O@     X�@     �l@     Ȉ@      u@     �@@      1@     @l@     t@      0@     �B@     Pt@      G@     w@     `h@     pw@      l@      9@      1@     �e@     �l@      .@     �@@     �o@      C@     �j@     �a@      q@      f@      7@      �?      H@     �R@      �?       @      Q@      @     @Y@      =@     @X@     �@@      �?      �?      :@      <@              �?      H@       @      I@      (@      O@      2@      �?              6@      G@      �?      @      4@      @     �I@      1@     �A@      .@              0@     @_@     �c@      ,@      9@      g@     �@@      \@      \@     �e@     �a@      6@      @     �W@     �`@      "@      7@     �a@      6@     �X@     �S@      c@     �W@      0@      $@      ?@      7@      @       @     �E@      &@      ,@     �@@      6@     �H@      @             �J@     �V@      �?      @      R@       @     �c@      K@     �Y@      H@       @              .@      2@                      *@      @     �P@      @     �C@      *@      �?              ,@      0@                      *@      �?     �J@              A@      &@                      �?       @                              @      *@      @      @       @      �?              C@      R@      �?      @     �M@      @     �V@     �I@      P@     �A@      �?              &@      F@      �?      @      5@              P@      :@     �C@      0@                      ;@      <@                      C@      @      :@      9@      9@      3@      �?              [@     �l@      @      .@     �c@      0@     Ѓ@     �A@      z@      \@       @             @R@     �f@      @      "@      X@      ,@     h�@      0@     �s@     @Q@      @              ;@      J@                      2@      $@     �W@      @     �L@      ,@      @              $@      :@                      2@      @     @P@      �?      H@      $@                      1@      :@                              @      >@      @      "@      @      @              G@     ``@      @      "@     �S@      @     �|@      &@     0p@     �K@      �?              :@     �Q@       @              @@             Pt@      @      e@      ;@                      4@      N@      @      "@      G@      @      a@      @     �V@      <@      �?             �A@      G@              @      N@       @     @S@      3@     �Y@     �E@      @             �@@      F@              @     �G@       @      K@      ,@     @U@      D@      @              5@      B@              @      <@      �?     �C@      ,@     @S@      >@      @              (@       @                      3@      �?      .@               @      $@                       @       @               @      *@              7@      @      1@      @                              �?                      @              .@              $@      �?                       @      �?               @      @               @      @      @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJCp{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?n'��8@�	           ��@       	                    �?�I9H	@           T�@                           �?�9�I@-           0~@                          �6@#�JO�@s            �g@������������������������       ��!2�T@?            �X@������������������������       �j|=�J@4             W@                          �6@
�Q"v�@�            @r@������������������������       �)i#�@k            �d@������������������������       �y�q�s@O             `@
                          �4@}��E�	@�           ȑ@                          �3@��f�B�@           �y@������������������������       �pM��C�@�            `s@������������������������       �f�{��@?            @Y@                           �?�S��	@�           ��@������������������������       �+��"@-             Q@������������������������       �]�
�	@�           ��@                          �5@�@*�-�@�           �@                          �4@����8@y           @�@                           @Pf�i�@�           ��@������������������������       ����R�@=           ��@������������������������       ��I-R�� @�           0�@                            �?]�J�@�            `j@������������������������       ��=��G@N             ]@������������������������       ��	m7��@6            �W@                           @����+g@            �@                          �=@��Ȧ@�             o@������������������������       �7�B{Re@�            @k@������������������������       �NQTd��@             >@                           @~�����@�           `�@������������������������       �&����U@�            �y@������������������������       ���_1v@�            `j@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �s@     ��@      <@      P@     �}@     �P@     x�@     `l@     H�@     u@      :@      0@      f@     �o@      7@     �E@     �n@     �C@      k@      b@     `p@     �f@      6@      �?     �I@     @R@      @      &@     �N@      �?     �Z@      A@     �V@      I@       @      �?      6@      8@                      :@              K@      $@     �B@      0@      �?               @      $@                      @              D@      @      :@       @              �?      4@      ,@                      3@              ,@      @      &@       @      �?              =@     �H@      @      &@     �A@      �?      J@      8@     �J@      A@      �?              1@      7@       @      @      1@              H@      "@      8@      2@      �?              (@      :@      �?      @      2@      �?      @      .@      =@      0@              .@     @_@     �f@      4@      @@     �f@      C@     �[@     �[@     �e@     �`@      4@      @     �@@      E@      @       @     @R@      @     �K@     �C@     @V@     �I@      @      @      7@      A@      @      @     �H@      @     �F@      >@      N@     �G@       @              $@       @      �?       @      8@              $@      "@      =@      @      @      $@      W@     `a@      0@      8@     �[@      @@     �K@     �Q@     �T@     @T@      ,@      @      .@      @              @      4@      @      �?      @      @       @              @     @S@     �`@      0@      5@     �V@      9@      K@     @P@     �S@     �S@      ,@             �a@     r@      @      5@     �l@      ;@     ��@     �T@     �@     `c@      @             �O@     �g@      @      *@      ]@      $@     p�@      @@      w@     @Q@      @              O@     @b@      @      (@      V@      @     �@      <@     �r@      O@                      E@      R@       @      @      I@      @      g@      4@     �^@      @@                      4@     �R@      �?      @      C@              t@       @     �f@      >@                      �?      E@              �?      <@      @      J@      @     �P@      @      @              �?      ;@              �?      @      @      ?@      @     �B@       @      �?                      .@                      5@      �?      5@              =@      @      @             �S@     @Y@       @       @      \@      1@      m@     �I@     `f@     �U@                     �E@      3@                     �A@      @     �J@      :@     �E@      6@                     �C@      0@                      ?@      @      G@      2@      E@      5@                      @      @                      @       @      @       @      �?      �?                      B@     �T@       @       @     @S@      $@     �f@      9@      a@      P@                      5@      L@              �?     �H@       @     �a@      0@     @T@      D@                      .@      :@       @      @      <@       @     �B@      "@     �K@      8@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJY�.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @]L*�X@�	           ��@       	                    �?��S���@v           �@                           �?e�w+S@�           ��@                            �?�ʤ�@�            �t@������������������������       ��q{��@<            @\@������������������������       ��d��ڟ@�             k@                            �?�ex�k@�            @u@������������������������       �F���@s            �g@������������������������       ��].�@`            �b@
                          �8@��B~	@�           ��@                          �2@���%	@�            �@������������������������       ���@K@�            �r@������������������������       ��s�e	@�           ��@                            �?��Ǽ��	@           �z@������������������������       ���f�/�@�            @l@������������������������       ���w7�E
@�             i@                           �?�F*"3@=           �@                          �4@
-��� @r           ȁ@                           �?��Te��?�            @u@������������������������       �����݀�?�            �i@������������������������       �A+�4Պ�?]             a@                          �5@� �@�            �l@������������������������       �m�-}ݚ�?#            �K@������������������������       ��Ղ�v@l            �e@                            �?x�w��@�            �@                           @J��i@�           p�@������������������������       ����.��@�           ��@������������������������       ��swn`P@	             .@                           @���
,�@A           �@������������������������       ���Y��B@�            �w@������������������������       �� +	Vc@U             `@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     p�@      9@      H@     �|@     �U@     `�@     @m@     ��@     w@      B@      2@     �i@     �s@      3@      @@      t@     �O@     @w@     �h@     0v@     `o@     �@@      �?      L@     �U@       @      @     �S@       @     �e@      A@     @c@     @Q@      �?      �?      :@     �C@       @      @     �D@      @     �V@      3@     �P@      ?@              �?      @      5@              @      .@      @      A@       @      6@      @                      6@      2@       @      @      :@      �?     �L@      1@     �F@      9@                      >@      H@                      C@       @     @T@      .@     �U@      C@      �?              1@      >@                      &@              D@      @     �P@      3@      �?              *@      2@                      ;@       @     �D@      &@      4@      3@              1@     �b@      m@      1@      9@      n@     �K@      i@     @d@      i@     �f@      @@       @     �]@     �d@      &@      1@     �g@      >@     `e@      X@      c@     �[@      6@       @      8@      F@       @              E@      @     @Q@     �@@     �I@      ?@      �?      @     �W@     @^@      "@      1@     @b@      ;@     �Y@     �O@     @Y@     �S@      5@      "@      @@     �P@      @       @     �J@      9@      =@     �P@     �H@      R@      $@       @      2@      >@      @      @      @@      $@      *@     �D@      =@     �D@      �?      @      ,@     �B@      @       @      5@      .@      0@      9@      4@      ?@      "@             @T@     �m@      @      0@     �a@      8@     ��@      C@     �z@     �]@      @              .@     �T@              @      6@      @     �q@      "@     @^@      <@                      &@      D@              @      "@             �g@      @     �Q@      $@                      @      5@              @      @              \@       @      F@       @                      @      3@                      @             �S@       @      :@       @                      @     �E@                      *@      @     �V@      @     �I@      2@                              3@                      @              2@      �?      &@                              @      8@                      @      @     @R@      @      D@      2@                     �P@     �c@      @      &@      ^@      4@     �u@      =@     Ps@     �V@      @              C@     @T@              @      N@      *@      j@      .@     �f@     �J@                     �B@     @T@              @      N@      @     �i@      *@     @f@     �J@                      �?                       @              @      �?       @      @                              <@     �R@      @      @      N@      @     �a@      ,@      `@     �B@      @              6@     �M@              @     �E@       @     �]@      $@     �X@      5@      �?              @      0@      @      @      1@      @      8@      @      =@      0@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��6hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �??��w�t@�	           ��@       	                    �?�#f�s	@           T�@                           �?N-{�@4           �~@                           �?�s�{�@z             h@������������������������       �N�=�O@4            �T@������������������������       ��;T�u�@F            @[@                            �?:'�C
�@�            �r@������������������������       ����e��@`            �c@������������������������       ����s�@Z            �a@
                           �?tV��1
@�           ��@                          �=@��%�PM@
            z@������������������������       ����!@�            Px@������������������������       ���V)}�@             =@                          �7@��k0�
@�           @�@������������������������       ���s  
@�             x@������������������������       ���e��
@�            �t@                          �2@���!{@�           �@                           �?!?���@�           ��@                          �1@��sg|@�            �v@������������������������       ��¢��L@�            �n@������������������������       ���L�@J            @\@                           �?O��1�@�            �v@������������������������       �z*w��?O             `@������������������������       ��?�d)
@�            @m@                           @�D$�@�           ��@                          �>@JTƮ��@	           �y@������������������������       ��b�n�@�            `x@������������������������       �_��˂ @             4@                            �?�V_��V@�            �@������������������������       �@Zu��@�           x�@������������������������       �l�U��@K           Ȁ@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     ��@     �@@      M@      }@      S@     �@      m@     ��@     �u@      D@      4@     �e@      m@      5@      B@      n@      F@     `l@     �b@     �p@     �e@      @@      �?     �H@     �R@      @      @     @Q@      �?     �Z@      =@     @Z@      F@      @      �?      $@      >@                      ;@             �H@       @      J@      .@              �?       @      (@                      *@              9@      @      8@      @                       @      2@                      ,@              8@      @      <@      (@                     �C@      F@      @      @      E@      �?      M@      5@     �J@      =@      @              1@      6@              @      2@              9@      .@     �@@      2@      @              6@      6@      @      �?      8@      �?     �@@      @      4@      &@              3@     �_@     �c@      2@      ?@     `e@     �E@      ^@      ^@     �d@     @`@      <@      �?      =@     @R@       @      $@     �R@       @     �L@      E@     @P@      J@      @      �?      :@     @R@       @      $@     �Q@      @     �K@      A@      O@      F@      @              @                              @       @       @       @      @       @              2@     @X@     �U@      0@      5@     @X@     �A@     �O@     �S@      Y@     �S@      7@      &@     �L@     �L@      "@      &@     �K@      @      E@      A@      L@     �B@       @      @      D@      =@      @      $@      E@      <@      5@      F@      F@     �D@      .@             @_@     �r@      (@      6@      l@      @@     Ї@     �T@     8�@      f@       @              5@     �T@      �?      @     �B@             �t@      3@     �d@     �I@      @              (@     �E@              @      <@             �c@      (@     �S@      :@                      @      B@              @      0@              \@      &@     �H@      *@                      @      @                      (@              G@      �?      =@      *@                      "@      D@      �?       @      "@              f@      @     @V@      9@      @              @      @                      @             �R@              8@       @      @               @     �@@      �?       @      @             �Y@      @     @P@      1@                      Z@     �j@      &@      1@     `g@      @@     �z@      P@      x@     �_@      @             �A@      O@       @      @      J@      &@     @V@     �@@     @R@     �G@      �?             �A@      M@       @      @      G@      &@     �T@      ?@     @R@     �G@      �?                      @              �?      @              @       @                                     @Q@     �b@      "@      (@     �`@      5@     0u@      ?@     ps@     �S@      @              E@      U@      @       @     �R@      ,@     �d@      7@     `d@      H@      @              ;@     �P@      @      $@     �N@      @     �e@       @     �b@      ?@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���c@�	           ��@       	                   �2@�<)���@           ��@                          �1@��&	q @           p{@                            @�Hd/N7�?�            �p@������������������������       ��Io=�?�             k@������������������������       ��8t�;�?$            �J@                           @��`y��@h             e@������������������������       ���4��c@5            @T@������������������������       ���;w�7�?3             V@
                          �<@��V-�@           ��@                          �3@�R�@�           ��@������������������������       ��>�-��@P            �^@������������������������       ��n�7@r           Ђ@                          �>@�w��@?            @W@������������������������       ���B�o�@"            �J@������������������������       �mg��1@             D@                           @�A��,*@�           ¤@                          �5@TF�)@�           ��@                           �?�$8S<�@           ؓ@������������������������       ��ʢY�@$            }@������������������������       �I��ݶ�@�           0�@                          @@@����i!	@�           H�@������������������������       �z���@�           ��@������������������������       �>��F�@@             C@                          �3@�}x�@�            �q@                          �1@h!{w�@,            �R@������������������������       ��m@             9@������������������������       �ǀd�F&@             I@                            @r���S7@�            �i@������������������������       � ��
r@l            �c@������������������������       �w�dk�@!            �H@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     Pp@     h�@     �@@     �J@     @|@     �U@     l�@      h@     (�@     �w@      @@             @S@     `e@       @      "@     @Y@       @     P~@      B@     �r@      O@      @              ,@      I@              �?      6@      �?     �l@      &@      W@      2@                      "@      A@              �?      ,@              c@      @     �I@      @                       @      >@              �?      *@             @^@      �?      D@      @                      �?      @                      �?              @@       @      &@       @                      @      0@                       @      �?     @S@       @     �D@      *@                      @       @                      @      �?      6@      @      9@      $@                      �?       @                      �?             �K@      @      0@      @                     �O@     @^@       @       @     �S@      @     �o@      9@      j@      F@      @             �K@     �Z@       @      @     �Q@      @     �m@      .@     `h@      :@       @              @      ,@                      @      �?      @@      @     �J@      @                     �H@     @W@       @      @     @P@      @     �i@      $@     �a@      4@       @               @      ,@              �?      "@      �?      0@      $@      ,@      2@       @              @      (@                      @              &@      @      $@      "@       @              @       @              �?      @      �?      @      @      @      "@              (@      g@      x@      ?@      F@     �u@     �S@     ��@     �c@     �@     �s@      <@      (@     `c@     �u@      ?@      F@     �s@     @P@     �@     �`@     `}@     `q@      3@       @     �M@     �h@      1@      3@      a@      7@     �u@      Q@     pq@     �]@       @       @     �A@      M@      "@      0@     �S@      &@     �Q@      G@      Q@      Q@       @              8@     �a@       @      @     �M@      (@     0q@      6@     `j@     �I@              $@      X@     �b@      ,@      9@      f@      E@     @d@     �P@     �g@     �c@      1@      @     �V@     `b@      (@      9@     �e@      A@      d@     @P@     �g@     @b@      1@      @      @      �?       @              @       @      �?      �?              *@                      =@     �C@                      C@      ,@      M@      6@      A@      C@      "@              @      @                      "@      @      9@       @      @      1@      @              @                               @      @      @      �?      @      @                              @                      @       @      4@      �?      �?      &@      @              :@      A@                      =@      "@     �@@      4@      <@      5@      @              4@      7@                      6@      @      9@      1@      4@      5@      @              @      &@                      @      @       @      @       @               @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ!�<PhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��Q�$w@�	           ��@       	                    �?�m�p&	@s           0�@                          �<@a�\Y�@�           �@                           �?-� Il@s           x�@������������������������       ���C�@�             q@������������������������       �]/2UWy@�            �s@                          @@@]���@0            �S@������������������������       ��MP���@&             P@������������������������       ���Z-�@
             ,@
                          �3@��WȪ	@�           �@                           �?�_��QK@           �|@������������������������       �-*(�	@�            ps@������������������������       �j?��e@`            �b@                           @��1�	@�           ��@������������������������       �t�zٹ�	@T           ��@������������������������       �)DH �	@c            �c@                           �?u
���@D           Ě@                          �4@M= � @j           0�@                           @���aϭ�?�            �u@������������������������       �
�Z���?�            `o@������������������������       �f�F��_@?            �X@                           �?��[�-�@�             i@������������������������       ��₲C@N            @\@������������������������       �xg��@8            �U@                           @˒�:@�           ,�@                          �7@
bp�b@            �@������������������������       �Zை�g@�           �@������������������������       �e��bB@}            `h@                            �?�Vҿ%�@�            �t@������������������������       �@!	B@1            �T@������������������������       ���/U�@�             o@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      r@     0�@      ;@      O@      {@     �W@     ��@     �m@     ��@     �v@      B@      1@     `i@      t@      3@      H@     �r@     �R@     �v@     �g@     �w@      o@     �@@      �?      M@     @W@       @      &@     �Q@      @     �c@     �B@     �c@     �Q@      @      �?     �H@     �U@       @      @      O@      @     �c@      9@      b@     �H@      @      �?      9@     �D@       @      @      A@      @     �T@      2@      E@      0@       @              8@     �F@               @      <@             @R@      @     �Y@     �@@       @              "@      @              @      "@              @      (@      (@      5@      �?              @      @                      @              @      $@      (@      5@      �?               @       @              @      @                       @                              0@      b@     �l@      1@     �B@     �l@     �Q@     �i@     �b@      l@     `f@      <@      @      9@      R@      �?      $@     �P@      &@      Y@      G@     �P@      J@      @      @      4@      E@      �?       @      J@      $@      L@      ?@     �D@     �C@      @              @      >@               @      ,@      �?      F@      .@      9@      *@              (@      ^@     �c@      0@      ;@     `d@     �M@     @Z@     @Z@     �c@     �_@      5@      @     �X@     �a@      0@      9@      a@      J@     �V@     @Q@     �b@     �[@      0@      @      5@      .@               @      :@      @      .@      B@       @      1@      @             @U@     �l@       @      ,@     �`@      3@     P�@     �H@     �{@     @\@      @              4@     �R@              �?      8@      @      q@      "@      _@      4@      �?              ,@      H@              �?       @             �g@      @     �Q@      (@      �?              "@      ?@                      @             �b@       @     �H@      @                      @      1@              �?      @             �C@      @      6@      @      �?              @      :@                      0@      @     �U@       @     �J@       @                      @      (@                      &@       @     �I@      �?      =@       @                      �?      ,@                      @      �?     �A@      �?      8@      @                     @P@     @c@       @      *@     �[@      0@     �u@      D@     �s@     @W@       @             �E@     �Z@      @      @     �Q@       @     0r@      5@      k@      Q@       @              <@      U@      @       @     �C@       @     �m@      (@     @e@     �I@      �?              .@      6@              �?      @@              J@      "@      G@      1@      �?              6@      H@      @      $@     �C@       @     �J@      3@     �Y@      9@                      "@      &@              �?      @      �?      4@       @      8@      @                      *@     �B@      @      "@      B@      @     �@@      &@     �S@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ^AFghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @G��|--@�	           ��@       	                   �3@�,%�տ@`           ��@                          �1@���@�           �@                            �?W�nx@�            `n@������������������������       ��5�Ie@3            �U@������������������������       ���e��@m            �c@                           �?�;��d�@�            �x@������������������������       �#ۘ30>@V            @a@������������������������       ������@�            @p@
                            @A�G
5	@�           x�@                           �?E��<	@H           �@������������������������       �G�x��@�            �o@������������������������       �В�5�	@�            �@                          �=@b��%�@�           ��@������������������������       �f��K�@V           ��@������������������������       ������	@+             O@                           @'o��@T           ��@                          �4@��H�<�@�           ��@                           �?1?!} @�           `�@������������������������       �F\�ֆ��?�             p@������������������������       �Q8��@           �|@                          �8@I��.��@C            @������������������������       �%�;�mz@�            `s@������������������������       ���8��q@{            �g@                           �?��~��#@W           `�@                            @�|���@�            Pr@������������������������       ��!��@�            @j@������������������������       �U$O �@,            �T@                          �7@_+��fJ@�            pp@������������������������       �o�5Ԛf@t            �f@������������������������       ����*@5             T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     @r@     ��@      9@      H@     `}@     �V@     P�@     �h@     ȉ@     `w@      9@      3@     @i@     �s@      0@     �C@     �s@     �R@     `u@      c@     �x@     @o@      5@      @      J@     @X@              @     �R@      0@     @b@      D@     �^@     @U@              @      0@      E@              �?      5@      �?     @R@      (@     �H@      9@                      @      2@                      �?      �?      ;@      �?      5@      &@              @      "@      8@              �?      4@              G@      &@      <@      ,@              �?      B@     �K@              @     �J@      .@     @R@      <@     @R@      N@                      .@      7@              �?      "@      �?      =@      @      C@      2@              �?      5@      @@              @      F@      ,@      F@      8@     �A@      E@              .@     �b@     `k@      0@      A@     �n@     �M@     �h@      \@     �p@     �d@      5@       @      V@      ]@      @      7@     �b@      I@     �^@     �P@     `c@      Z@      &@              =@     �B@              @      ?@      @     �M@      $@      M@      4@      �?       @     �M@     �S@      @      3@     �]@     �F@      P@      L@     @X@      U@      $@      @      O@     �Y@      &@      &@      X@      "@     @R@      G@     �\@     �N@      $@      @      M@     �U@      $@      @     �U@      @     �P@     �E@     �[@     �J@      $@      @      @      0@      �?      @      "@       @      @      @      @       @               @     �V@     `l@      "@      "@     �b@      .@     ��@      G@     {@      _@      @       @      H@     `d@       @       @     �V@      $@     `@      9@     �r@     @P@       @              8@     @X@       @      �?      >@              v@      $@      e@      ?@                      @      =@                       @             `d@      @      F@      @                      4@      Q@       @      �?      6@             �g@      @     @_@      ;@               @      8@     �P@              �?      N@      $@     �b@      .@     �`@      A@       @       @      .@     �H@                      B@      "@     �Z@      @     �Q@      1@       @              "@      1@              �?      8@      �?      F@      &@      P@      1@                      E@      P@      @      @     �N@      @     �c@      5@     @`@     �M@       @              6@     �@@      @      @     �B@      �?     @W@      @      M@      @@                      4@      =@       @      @     �A@             �K@      @     �F@      0@                       @      @      @       @       @      �?      C@       @      *@      0@                      4@      ?@       @       @      8@      @     @P@      ,@      R@      ;@       @              ,@      9@              �?      2@      @     �L@      @     �E@      ,@       @              @      @       @      �?      @      �?       @       @      =@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�>�OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�A��L@�	           ��@       	                   �;@?����@Y           d�@                           �?��Yl��@�           ؝@                          �5@-�*�\@J           ��@������������������������       �u#}��@�           ��@������������������������       ��d朅@s           x�@                           �?��+�#t@E           ��@������������������������       �E��-�U@U            `a@������������������������       �E#5@��@�            Px@
                           �?T�G�
@�            �s@                          �<@����	@K             \@������������������������       ����VC@             B@������������������������       �b�)R@4             S@                          �<@`�us�N
@            �i@������������������������       �q(||@
@             G@������������������������       ��X�LJ	@e            �c@                           @���j#@?           \�@                          �7@��;��@*           ��@                           �?�a��A@3           ��@������������������������       � �O�=��?'           �{@������������������������       �S�ꅮ.@           �@                           �?��`v�@�            �x@������������������������       ��GbY�S@|            �j@������������������������       �UKZf��@{             g@                           �?I���Y�@             D@������������������������       �>��_� @             0@������������������������       ��T�}
@             8@�t�bh�h5h8K ��h:��R�(KKKK��h��B 
        2@     �r@     �@      :@     �I@     @}@     �U@     P�@      k@     ��@     @w@      ?@      2@     �i@     `t@      5@     �A@      v@     �M@     @x@      f@     �v@     p@      8@       @      e@     �q@      .@      6@     �s@     �A@     �v@      b@     �t@      i@      3@       @     ``@     �i@      .@      1@     @o@      :@     �k@     �Y@     `m@     �b@      2@      @     �J@     �Z@      $@       @     @a@      (@     �b@     �J@      b@     �Y@      @      �?     �S@      Y@      @      "@      \@      ,@     �Q@      I@     �V@      H@      *@             �B@     �S@              @      Q@      "@     �a@      E@     �W@      I@      �?              *@      (@                      .@      �?      H@      �?     �B@      (@                      8@     �P@              @     �J@       @     �W@     �D@     �L@      C@      �?      $@     �C@      D@      @      *@      B@      8@      7@      @@      ?@     �L@      @       @      (@      4@      �?      @      3@      (@       @       @      @      3@              @      @      @      �?              &@      @      �?      �?      @       @              @      "@      ,@              @       @      "@      �?      @      �?      1@               @      ;@      4@      @       @      1@      (@      5@      8@      9@      C@      @       @      @      @      @       @       @       @      @              @       @      @              6@      *@       @      @      .@      $@      .@      8@      4@      >@      �?             �V@     �k@      @      0@     �\@      ;@     0�@      D@     `{@     �\@      @             �T@     �k@       @      .@     �Z@      2@     �@      B@     @{@     @\@      @              J@     �e@       @      @     �L@      $@     H�@      0@     �t@     �Q@      @              &@      J@               @      .@      �?     �m@      @     @X@      5@      �?             �D@     �^@       @      @      E@      "@     �q@      "@     �m@      I@      @              ?@     �F@              $@     �H@       @     �V@      4@     �Y@      E@      �?              8@      =@              @      0@      @     �L@      @      H@      7@      �?              @      0@              @     �@@      @     �@@      ,@     �K@      3@                      @      �?      @      �?       @      "@      @      @       @       @                                              �?       @       @      �?      @              �?                      @      �?      @              @      �?       @      �?       @      �?        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?/��I�F@�	           ��@       	                    �?N�ɳ�	@�           ��@                           �?���Q�@�           h�@                           �?*;d���@�            �o@������������������������       ���[ܕ@:             T@������������������������       ���V*!	@h            �e@                           �?�·��@�            �v@������������������������       ������a@<            �V@������������������������       ����W�j@�            @q@
                          �;@Z~�'�	@f           ��@                           �?�v�׎	@�            �@������������������������       �VE���^@�            �m@������������������������       ���晖�	@`           ��@                          �<@& ��O	@s            `f@������������������������       �Rga���@             C@������������������������       �4�(P`�@]            �a@                           �?Zက��@�           R�@                          �4@�DM�av@�           ��@                          �0@^P��EB @           �{@������������������������       ���Ѿz�?*            �P@������������������������       �e��ק� @�            �w@                            �?�{��@�            @t@������������������������       �w?�.�� @-            �S@������������������������       �Q�m �@�            �n@                           @$����@�           ��@                          �9@�%��&y@�           ��@������������������������       �B^6��@i           Ё@������������������������       ��wW*��@O            �`@                           @-hw�B@           h�@������������������������       ��G���"@K           �@������������������������       ����t@�            �t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �r@     h�@      :@     �M@     �z@     @Y@     ,�@     `f@     H�@     @v@     �D@      3@     `d@     `i@      *@     �B@     @l@     �P@     �k@     �]@     q@     �h@      @@       @     �I@     @T@      @      (@     �W@      3@     �^@      E@     �]@      O@       @       @      :@     �@@               @     �F@      &@     �H@      ,@     �B@      ;@      @      �?       @      @                       @              ?@      @      3@      @              @      2@      <@               @     �B@      &@      2@      $@      2@      7@      @              9@      H@      @      $@     �H@       @     @R@      <@     �T@     �A@      @              @      .@                      0@              1@      �?      <@      @      @              3@     �@@      @      $@     �@@       @      L@      ;@      K@      ?@       @      &@      \@     �^@      $@      9@     �`@     �G@     �X@     @S@     @c@     �`@      8@      @      V@      Z@      @      2@     @[@      >@     @U@      Q@     �a@     �V@      8@              5@      B@      @      @      B@             �E@      1@     �J@      6@      @      @     �P@      Q@       @      .@     @R@      >@      E@     �I@     �U@      Q@      3@      @      8@      2@      @      @      7@      1@      ,@      "@      ,@      F@               @       @      @       @              @      @       @              �?      $@               @      6@      *@      @      @      4@      (@      @      "@      *@      A@               @     �`@      t@      *@      6@     �i@     �A@     p�@      N@     ��@      d@      "@              9@     �X@       @       @      H@      @      v@      ,@     `h@      5@      @              0@     �G@               @      5@              l@      @     @[@      ,@       @                      ,@                                     �B@              (@      @                      0@     �@@               @      5@             �g@      @     @X@      &@       @              "@      J@       @              ;@      @     �_@       @     �U@      @       @                      ,@       @              @              A@      �?      4@               @              "@      C@                      5@      @     @W@      @     �P@      @               @     �[@     �k@      &@      4@     �c@      ?@     �|@      G@     Pw@     `a@      @       @      P@      \@      @      $@     @S@      :@     �d@     �@@     �a@     �P@      @       @     �G@      X@      @      @     �J@      3@      c@      8@      ]@      H@      @              1@      0@              @      8@      @      (@      "@      9@      2@                      G@     �[@      @      $@      T@      @     �r@      *@      m@     @R@       @              2@     �O@               @      H@             `k@      &@     @c@      ?@      �?              <@      H@      @       @      @@      @     �S@       @     �S@      E@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���yhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?����:@w	           ��@       	                     @��
ū�@�            �@                          �4@Oۍ�b�@%            �@                            �?#��u@/           �@������������������������       �T���c�?o            �h@������������������������       ���_)��@�            `s@                          �<@���'@�            �x@������������������������       �ѕ/���@�            �t@������������������������       �`��>� @(            @P@
                          �6@-���Q@�            �s@                          �2@�]'.=�@�            �i@������������������������       ���|
��?D             [@������������������������       �1�ܿ@@            �X@                           @:��b�@H            �[@������������������������       ���ߞ��@<            �V@������������������������       ��r?I���?             3@                          �4@{:�@�F@�           �@                          �1@���'h@�           ��@                           �?�$����@�            px@������������������������       �I��u�@s            `g@������������������������       �<͞�p@�            �i@                           @��[�\@           ��@������������������������       �#�[�@`           ��@������������������������       �2b~d�@�             o@                           @�O,u�R	@�           (�@                           �?���f�	@P           @�@������������������������       �6-���#@�            �p@������������������������       �cr��-
@�           ȅ@                           @S�L��@A           �@������������������������       �WC���@�            �u@������������������������       �%L{��@f            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �r@     ��@      B@     �N@     �z@     @S@     ��@     �h@     ��@     �t@     �C@             �U@     `c@      �?      $@     �Y@      $@     �~@      C@     `p@     �I@       @             �M@     �_@      �?      @     �P@      $@     pv@      ;@     �h@     �D@       @              6@      P@              �?      :@      �?      p@      "@     �Y@      3@      @              @      9@              �?      @             �Z@      @      F@      $@                      3@     �C@                      6@      �?      c@      @      M@      "@      @             �B@      O@      �?       @     �D@      "@     @Y@      2@     @X@      6@      @              ?@     �G@      �?      �?     �B@       @     @W@      &@     �V@      $@                      @      .@              �?      @      �?       @      @      @      (@      @              <@      =@              @     �A@             �`@      &@     �O@      $@                      8@      1@              @      *@             @Y@      @     �C@      @                      $@      @              �?      "@              O@       @      1@       @                      ,@      (@               @      @             �C@      �?      6@      @                      @      (@              @      6@              @@       @      8@      @                       @      (@              @      6@              3@      @      7@      @                       @                                              *@      @      �?                      2@     �j@     �y@     �A@     �I@      t@     �P@      �@      d@     P�@     �q@      ?@       @     �P@     �g@      &@      &@      ^@      3@     �u@     �M@     �p@     �\@      (@              3@      Q@      �?      �?      2@      �?      a@      *@     �W@     �C@                      "@      D@      �?      �?      @      �?     �R@      @      A@      0@                      $@      <@                      &@             �O@      "@      N@      7@               @     �G@     @^@      $@      $@     �Y@      2@     `j@      G@     @e@     �R@      (@      �?     �B@     �U@       @      @      U@      ,@      b@      4@     @^@     �I@              �?      $@      A@       @      @      2@      @     �P@      :@     �H@      8@      (@      0@     �b@     �k@      8@      D@     @i@      H@      m@     �Y@      p@     @e@      3@      0@     @\@      d@      1@      =@      `@      D@     �Z@      V@     �`@      _@      *@       @      &@     �F@      @      @     �C@      @      D@      5@     �E@     �J@      @      ,@     �Y@     �\@      ,@      6@     �V@      B@     �P@     �P@     �V@     �Q@      $@             �A@     �O@      @      &@     @R@       @     �_@      ,@     @_@      G@      @              <@     �C@      �?      @      J@      �?     �Z@      @     @T@      <@      �?              @      8@      @       @      5@      @      4@      @      F@      2@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�C�nhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �8@���ʖ@�	           ��@       	                    �?ȍ� �@m           2�@                          �5@�¡�<�@m           �@                            �?ǡ���@�           �@������������������������       �ܹ��|� @�             j@������������������������       �ϻi�ȅ@U           ��@                            �?5X<��@�            @k@������������������������       �� ���@M            �Z@������������������������       ����h@E            �[@
                           �?�����@            p�@                           �?؟�1H
	@Q            �`@������������������������       �2Z2x@             F@������������������������       �l5H��(	@6             V@                           @�z~F�A@�           `�@������������������������       ��Ԫ=��@           p�@������������������������       ����	@�            �o@                            �?HF�X��	@M           ��@                           �?:+X<	@8           8�@                          �;@j�'J��	@�            Pr@������������������������       �ۄk��@P            �`@������������������������       ��;��ya	@[             d@                           @�rc�>@�            @l@������������������������       �r�n�@y             h@������������������������       ��J�'�� @            �@@                          �=@E��>�	@           �z@                          �:@�.	@�            t@������������������������       ��2�6WG@k             e@������������������������       ��[B�@m             c@                          �?@����@=             Z@������������������������       �B�pn�@            �J@������������������������       ���S^�@            �I@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     ��@     �@@     �Q@     �z@      V@     ��@     �l@     ��@     u@     �A@      *@     `l@     �{@      1@     �H@     �r@     �I@     0�@      `@     ȃ@     �j@      3@             �P@     @a@       @      (@      P@      "@     �v@      7@     �l@     �F@      �?             �F@     �W@              &@      G@      "@     �s@      4@      e@      >@                       @      >@              �?      "@      @     @U@       @      Q@      "@                     �E@      P@              $@     �B@      @     �l@      2@     @Y@      5@                      6@      F@       @      �?      2@              I@      @      O@      .@      �?              ,@      &@      �?      �?      (@              :@      �?      @@       @      �?               @     �@@      �?              @              8@       @      >@      @              *@      d@     @s@      .@     �B@     �m@      E@     �@     �Z@      y@      e@      2@      @      *@      4@               @      :@      @      *@      (@      3@      *@                      @      &@                       @      �?      @              @      @              @       @      "@               @      2@      @      @      (@      ,@      @              "@     `b@      r@      .@      =@     �j@      C@     �~@     �W@     �w@     `c@      2@      @      _@     �n@      .@      9@     �f@      >@     �{@     �R@     �u@     �_@      $@      @      7@      F@              @      >@       @      H@      4@     �@@      =@       @      $@      S@     @b@      0@      6@     �_@     �B@     �]@      Y@      c@      _@      0@      @     �B@     �V@      @      $@      N@      5@      H@     �O@      V@      T@      $@      @      5@     �H@      @       @      D@      ,@      ,@      D@     �C@      H@      "@              $@      7@               @      ,@      "@      "@      =@      2@      (@      @      @      &@      :@      @      @      :@      @      @      &@      5@      B@      @              0@      E@               @      4@      @      A@      7@     �H@      @@      �?              $@      E@               @      3@      @      A@      (@     �E@      7@      �?              @                              �?                      &@      @      "@              @     �C@     �K@      $@      (@     �P@      0@     �Q@     �B@     @P@      F@      @       @      8@      B@      @       @     �G@      .@      N@      A@      M@      >@      @              *@      5@      @              8@      $@      7@      3@      D@      (@       @       @      &@      .@       @       @      7@      @     �B@      .@      2@      2@      @      @      .@      3@      @      $@      3@      �?      $@      @      @      ,@                      @      ,@      �?      @      ,@      �?      @      @      �?      @              @      &@      @       @      @      @              @              @      $@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJd[�ihG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?
�{|X@�	           ��@       	                    �?aJO;+�	@            �@                          �9@u��(�@�           �@                            �?�Ń�@3           �{@������������������������       ��R�M@]             a@������������������������       �$��w @�            Ps@                            �?"�F��n@R            ``@������������������������       �~�\9L>@             =@������������������������       ������@>            �Y@
                           �?���p
@�           Џ@                          �7@���{�
@�            `w@������������������������       �?=�~�@�            �k@������������������������       �;���+B
@f             c@                          �<@^�b
��	@�            �@������������������������       ���?sC�	@k            �@������������������������       ��F2�b@<             X@                          �4@_����@�           �@                           @�4��kw@           T�@                          �3@M���Lg@=           �~@������������������������       �U��㘀@�            �x@������������������������       �a�dO�W@A            �X@                            �?�׈Eڪ @�           H�@������������������������       ��Q��E� @�            y@������������������������       ����(�2 @�            �u@                          �7@������@�           �@                           �?�4\�S�@D           (�@������������������������       ��NTS�t@�            p@������������������������       ���zP�@�            @p@                           @��&o��@d           ��@������������������������       ���b�m@Q           x�@������������������������       �� J�G#@            �B@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     `�@      ?@     �K@      |@      V@      �@     �j@     ��@      u@      A@      6@     �e@     �j@      <@      ?@     �n@      I@     �l@     �a@     �o@     �g@      8@       @      C@      S@       @      "@      V@      0@      ]@      E@     �]@     �P@      @              @@      P@       @      "@     �Q@       @      X@      =@     �Y@      ?@       @              &@      3@              @      (@      @     �A@      @     �B@       @      �?              5@     �F@       @      @      M@      @     �N@      6@     �P@      7@      �?       @      @      (@                      2@       @      4@      *@      0@     �A@      �?      �?              @                       @      �?      @      @      @      �?              �?      @      "@                      $@      @      .@      "@      $@      A@      �?      4@     �`@      a@      :@      6@     �c@      A@     @\@     �X@     �`@     @_@      5@      @     �H@      O@      ,@      @      A@      0@      G@     �A@     �E@     �L@      @      @      ?@     �D@      @      �?      3@      @      E@      .@      =@      ;@      @      @      2@      5@      "@      @      .@      &@      @      4@      ,@      >@      @      *@     @U@     �R@      (@      1@     �^@      2@     �P@     �O@     �V@      Q@      .@      (@     @Q@     @P@      &@      "@      [@      *@     �O@      J@     @V@      F@      *@      �?      0@      "@      �?       @      ,@      @      @      &@      �?      8@       @             ``@     �u@      @      8@     �i@      C@     �@     @R@     ؀@     `b@      $@              H@     �g@      �?      @     �S@      @     ��@      :@     �q@     �O@      @              4@     �V@      �?      @     �C@      @     �e@      5@     @Y@     �B@                      1@      Q@              �?      1@      @     �b@      .@     @U@      @@                      @      6@      �?       @      6@              6@      @      0@      @                      <@     �X@              @      D@             �v@      @     �f@      :@      @              0@      J@              @      <@             �f@      �?     @Z@      (@                      (@     �G@                      (@              f@      @     �R@      ,@      @             �T@     `c@       @      1@     �_@      ?@     �p@     �G@      p@      U@      @              C@     �U@      �?      $@      I@      5@     @c@      @     �\@      ?@      @              5@      ?@              "@      <@      0@      U@      @     �F@      1@      @              1@     �K@      �?      �?      6@      @     �Q@      @     �Q@      ,@       @             �F@     @Q@      �?      @     @S@      $@      ]@     �D@     �a@     �J@       @              A@     �P@      �?      @     �P@       @      ]@     �@@     �a@     �J@       @              &@       @                      &@       @               @      @                �t�bub�     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJx>�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�*��/@�	           ��@       	                    �?	��3��@~           P�@                          �9@��n	z�@           �@                            @�R�в�@�           ��@������������������������       ��!�S^�@�             x@������������������������       �y@)υ�@�            �n@                           �?:�ӝ2>	@�            `i@������������������������       �[GI�;@@&             N@������������������������       ��� �WU	@Z            �a@
                            �?�Td�v@o           ��@                          �5@ȁ��X@�           x�@������������������������       �X���w�@�            �x@������������������������       ��Uv#�	@�            0v@                           @"�)vM@�           ��@������������������������       ��쓳��@r           ��@������������������������       �*�bW��@            �M@                           @qI��,@.           ��@                          �4@yD8{@�           ��@                           �?��.1A@�           p�@������������������������       ��@'�?�?�            `o@������������������������       �1"�h�[@	           0y@                            @�ij�"�@6           @������������������������       �%��I�@           �z@������������������������       �3?��)�?(             Q@                           @���;P�@W           �@                           �?V0��RU@�            0x@������������������������       �&���{ @�            �j@������������������������       ���l�G@k            �e@                            �?�j^��@j            �c@������������������������       ��c�6�R@6             U@������������������������       �#���Yz@4            �R@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �p@     `�@      ?@     �G@     @}@     @V@     ��@     `l@     ��@     �u@      ;@      .@     �g@     Pu@      6@      A@      t@      S@     �w@      g@     �x@      n@      4@      @      S@      _@      *@      @     @_@      A@      b@      S@     @]@      [@      @      @     �O@     �V@      @      �?     �Y@      .@      `@      M@     �W@     @P@      @      �?     �C@     �N@              �?     �M@      "@     �R@      G@      H@     �D@      @      @      8@      =@      @             �E@      @     �J@      (@      G@      8@      �?       @      *@      A@      @      @      7@      3@      0@      2@      7@     �E@                      @      *@               @      @              @      @      .@      ,@               @      "@      5@      @      @      4@      3@      $@      .@       @      =@              "@     @\@      k@      "@      <@     `h@      E@      m@      [@     �q@     �`@      .@      @     �O@      [@      @      3@     @S@      8@     �`@     �M@     �e@     �S@      @      �?      ;@     �F@       @      @      G@       @      W@      6@     �[@      B@      �?      @      B@     �O@      @      *@      ?@      0@      E@     �B@     �O@      E@      @      @      I@     @[@      @      "@     �]@      2@     �X@     �H@     �Z@     �K@      $@      @      F@     @V@      @      "@     @[@      ,@     @W@     �F@     @Z@      K@      @      �?      @      4@                      "@      @      @      @       @      �?      @             �R@     �n@      "@      *@     �b@      *@     �@     �E@     {@      Z@      @             �G@      g@                     �W@      "@     �z@      ;@     �r@      M@      @              6@      Y@                      @@      @      r@      *@     �d@      <@                      (@      ?@                      @             �a@      �?     �J@      @                      $@     @Q@                      9@      @     �b@      (@     @\@      6@                      9@      U@                      O@      @      a@      ,@     �`@      >@      @              9@     �T@                     �H@      @     �Z@      ,@     �\@      <@      @                      �?                      *@              >@              4@       @       @              <@     �O@      "@      *@      K@      @     `f@      0@     �`@      G@       @              0@      J@      "@      @      8@      �?      b@      (@     �W@      =@      �?              @      :@      @      �?      .@             �W@      @      I@      ,@      �?              *@      :@      @      @      "@      �?     �H@       @      F@      .@                      (@      &@               @      >@      @     �A@      @      C@      1@      �?               @      @              @      ,@      @      *@      @      ;@      @                      @       @              �?      0@              6@              &@      (@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ'<�OhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @}�+U��@�	           ��@       	                    �?��֐�@^           ^�@                           �?�)���b@�           ��@                          �<@ً<��,@*           0}@������������������������       ��氞�@           z@������������������������       ��s�t@"             I@                            �?�B��!@w            �g@������������������������       ��"�^VQ@+            �N@������������������������       ��CQ��@L             `@
                           @��{52s	@�           |�@                          �4@�˃Djd	@G           ��@������������������������       ��r����@O           @�@������������������������       �7�?�	@�           �@                           @K��!o@v            �f@������������������������       ��2��@�@T            ``@������������������������       ����,��@"            �I@                           �?���Q�d@B           h�@                          �2@p�'�d@m           �@                           @���.��?�            �m@������������������������       ���J�p��?o            �e@������������������������       �7%�&t@*             O@                            @�L��in@�            ps@������������������������       ���X�5\@�             q@������������������������       ���u>� @            �C@                           !@ߞR �r@�           ܑ@                           @�X�R@�           ��@������������������������       � +tT@�           �@������������������������       �\3���>@�            �t@������������������������       �������?             *@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@     �r@      �@      >@     �O@     @}@     �T@     H�@     @l@     @�@     w@      @@      4@     �j@     `v@      5@      F@     �s@      N@     @v@     �g@     `w@     `n@      >@             �Q@     @Z@       @      "@     �P@      @      e@      A@     @b@     �F@      @              K@      T@       @       @     �G@       @     @Z@      >@     �V@      E@      @             �G@     �R@       @      @      C@       @     @Y@      7@     �U@      =@      @              @      @              �?      "@              @      @      @      *@                      0@      9@              �?      3@       @     �O@      @      L@      @                       @      "@              �?      @      �?      6@              3@      @                      ,@      0@                      .@      �?     �D@      @     �B@                      4@     �a@     �o@      3@     �A@     @o@      L@     �g@     @c@     �l@     �h@      7@      0@     @_@     �k@      3@     �A@     �j@     �I@     @e@     @]@     `j@     �g@      0@       @      B@      U@       @      "@     �Q@      @      ^@      J@     �X@      N@      @      ,@     @V@     `a@      &@      :@     �a@      F@      I@     @P@      \@      `@      (@      @      2@      >@                      B@      @      2@     �B@      1@      $@      @              ,@      <@                      :@      @      ,@      ;@       @      @      @      @      @       @                      $@              @      $@      "@      @      @             @V@     @k@      "@      3@      c@      6@     (�@      C@      y@     �_@       @              2@      R@              @     �@@      @     �p@      @      ^@      9@      �?              @      3@               @      @             @b@             �I@      @      �?              @      $@                      �?             �^@              B@      �?                       @      "@               @      @              7@              .@      @      �?              *@     �J@               @      ;@      @     �]@      @     @Q@      3@                      $@     �H@                      :@      @     �X@      @     �N@      3@                      @      @               @      �?              4@      �?       @                             �Q@     @b@      "@      .@     �]@      0@     �u@      A@     �q@     @Y@      �?              P@      b@      "@      .@     @]@      ,@     �u@      A@     �q@     @Y@      �?              D@     �Z@      @      @     @Q@      @     �q@      4@     �g@     @R@                      8@      C@      @      &@      H@       @     @P@      ,@     �V@      <@      �?              @      �?                       @       @                      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��SnhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�q�*g@�	           ��@       	                   �1@�����@W           �@                           �?�Aza�@�           p�@                           @�d@�v @�            �o@������������������������       �kjR�T�?�            �i@������������������������       ���V�a�@             H@                           �?���/Y@�             w@������������������������       �?�ѳO@M             \@������������������������       ���S�o�@�             p@
                           �?�).F�@�           �@                           @{�f ��@I           ��@������������������������       ��5�	�^@�            �q@������������������������       ��Go<*�?�            �o@                           @����ޔ@t           `�@������������������������       ���Y��@�           ؃@������������������������       ��2�/�@�            w@                           �?2^���@R           `�@                          �8@� !�r@&            ~@                           �?�q�t#�@�            �k@������������������������       �i�o��@:            �U@������������������������       ��"S��@O             a@                           �?�4Ų��@�            p@������������������������       ��q7Ԧ�@O            @^@������������������������       �kG.�J�@N             a@                           @Ν�n�=	@,           ��@                           �?��.L��	@           ��@������������������������       �k���	@�            `k@������������������������       ���n��	@}           �@                          �<@�~y/�<@%           �}@������������������������       �����@�            �x@������������������������       �g%���@-             T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     `r@     Ѐ@      7@     �N@     �~@     �T@     Ȏ@     @i@     �@     �w@     �B@      @     @]@     pr@      "@      9@     �k@      ?@     ȅ@     �V@      ~@      e@      0@      @      6@     �T@      �?      @     �I@      �?     @p@      ,@     `a@     �E@      �?              @      ?@               @      8@             �_@      @      J@      "@      �?              @      >@                      ,@              Z@       @     �G@      @                      �?      �?               @      $@              6@       @      @      @      �?      @      1@      J@      �?       @      ;@      �?     �`@      $@     �U@      A@              @      &@      *@      �?       @      ,@      �?      6@      @      ;@      .@                      @     �C@                      *@              \@      @      N@      3@              @     �W@     �j@       @      5@     �e@      >@     P{@     @S@     pu@     �_@      .@              >@      R@      @      @     �A@      @      k@      7@     �]@      :@                      9@     �A@      @      @      ;@      @     �S@      2@     @P@      6@                      @     �B@                       @       @     `a@      @      K@      @              @     @P@     �a@      @      2@      a@      7@     �k@      K@      l@      Y@      .@      @     �H@      [@      @      ,@     �W@      7@     @V@      G@     �^@     �Q@      ,@              0@      @@       @      @     �E@             ``@       @     �Y@      >@      �?      0@      f@     `n@      ,@      B@     �p@      J@      r@     �[@      t@      j@      5@              F@     �Q@              &@      M@      $@     �^@      &@     @Z@     �F@      @              7@     �C@                      7@             @R@      @     �H@      (@                      "@      2@                      *@              0@      @      5@      @                      ,@      5@                      $@             �L@              <@      @                      5@      @@              &@     �A@      $@     �H@      @      L@     �@@      @              "@      ,@               @      &@       @      <@      @      9@      5@                      (@      2@              @      8@       @      5@      @      ?@      (@      @      0@     �`@     �e@      ,@      9@      j@      E@     �d@      Y@     �j@     `d@      2@      ,@     �V@     �^@      *@      ,@     �_@      ?@     �Q@     �S@     �Z@     �[@      1@      �?      *@      =@      @      @     �E@       @      =@      .@     �E@     �@@      @      *@     �S@     �W@       @      &@     �T@      =@     �D@      P@      P@     �S@      ,@       @      E@     �H@      �?      &@     �T@      &@      X@      5@      [@      J@      �?       @     �@@     �C@              @     �N@      &@     @V@      5@     �W@     �B@      �?              "@      $@      �?      @      5@              @              *@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��EM8@�	           ��@       	                    �?L|��8�@\           �@                          �8@����RK@�           h�@                          �6@��-�@            @}@������������������������       ����e@�             x@������������������������       �+���@2            �T@                          �<@���@p             g@������������������������       ��K��w@E             ^@������������������������       ��.��O@+            @P@
                          �2@�@�lȁ	@�           �@                           @�����@�            �r@������������������������       �N7D�@�            �i@������������������������       ��l����@<            @W@                           �?S���;�	@           4�@������������������������       �n_&"5@G            �_@������������������������       �74Bї�	@�           8�@                          �4@	�;ϋ@R           �@                           �?�v�E��@f           ��@                            �?0��W�?�            `w@������������������������       ����n��?;             X@������������������������       ���fMk��?�            `q@                           �?qzm�p@y           �@������������������������       �:� ��B@�             s@������������������������       �k,�v�@�            �r@                            @/�a�@�           ��@                          �5@��#��,@�           X�@������������������������       �ϱF�y�@]             c@������������������������       ���ǘ@7           0}@                           �?�����'@X            �`@������������������������       �s(��'8�?             E@������������������������       ��Ud�@@            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@      s@     ��@      5@      L@     �z@     �P@     ��@     `l@     p�@     pv@      E@      1@     `k@     @t@      1@     �F@      s@     �J@     `v@     @h@     @w@     `n@      A@             @P@     @Z@      �?      @      Q@      @     �e@      C@     `a@      G@      @              F@     @R@      �?              D@      �?     �a@      6@     @]@      =@      �?              A@     �P@                      8@      �?     �]@      5@     @W@      :@      �?              $@      @      �?              0@              5@      �?      8@      @                      5@      @@              @      <@      @     �@@      0@      6@      1@      @              &@      9@              @      3@      @      <@      @      .@      @       @              $@      @              @      "@              @      &@      @      &@       @      1@     @c@     `k@      0@      C@     �m@     �G@      g@     �c@      m@     �h@      =@       @      3@     �G@              �?      H@      @      H@      H@      M@      9@      �?      �?      "@      ;@              �?     �C@             �@@     �A@      G@      0@              �?      $@      4@                      "@      @      .@      *@      (@      "@      �?      .@     �`@     �e@      0@     �B@     �g@      F@      a@      [@     �e@     �e@      <@      @      2@      3@              &@      8@       @      @      @      8@      *@              $@     @]@      c@      0@      :@     �d@      E@     �`@     @Y@     �b@     �c@      <@             �U@     �m@      @      &@     �^@      ,@     x�@     �@@     �{@      ]@       @             �F@      a@      �?      @      D@      @     �{@      (@     `l@      N@       @              &@     �D@              �?      &@             @j@             @U@      *@       @                       @                      �?             @R@              0@      @                      &@     �C@              �?      $@              a@             @Q@      "@       @              A@     �W@      �?      @      =@      @      m@      (@     �a@     �G@                      2@     �E@      �?      @      3@              Z@      $@     @S@      <@                      0@      J@                      $@      @      `@       @     @P@      3@                      E@     �Y@      @      @     �T@       @     �j@      5@     �j@      L@      @              C@      X@       @      @     �R@      @     �d@      2@     @e@      E@      @              �?      <@                      3@       @      F@              J@       @      @             �B@      Q@       @      @     �K@      @     @^@      2@     �]@      D@                      @      @      �?      �?       @      �?     �G@      @     �F@      ,@       @                      �?                                      ;@       @      (@                              @      @      �?      �?       @      �?      4@      �?     �@@      ,@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�I�ghG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             @徆��b@�	           ��@       	                   �3@9A��S
	@x           ��@                           @G��]K@�           ��@                            @��ə�@(           �{@������������������������       ��<��F@�             q@������������������������       �� 0�R�@j            @e@                           @J6-,b@�             p@������������������������       �4��Y@>            @[@������������������������       �Q���bf@^            `b@
                           �?&��v�	@�           �@                            �?����01@           �x@������������������������       ��o.O@�            @k@������������������������       �f�:im@r            �e@                          �8@�����	@�           �@������������������������       ���X��C	@�           Є@������������������������       ����
f
@           z@                           @���gJ�@=           (�@                           @�oK)�x@�           ��@                           @2����%@�           L�@������������������������       �Ɖ��R�@           pz@������������������������       �A�
@�� @�           `�@������������������������       �p��E�"@             5@                            �?�X;�@[           �@                           �?�N��s}@K            �_@������������������������       ���� �?             J@������������������������       �&���n#@.            �R@                          �4@ybGq�@           @z@������������������������       ���vp"}@�            �g@������������������������       �uG�8�+@�             m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@      t@     ��@      @@     �P@     @{@      Q@     X�@     �l@     ��@     pu@     �A@      0@     �k@      t@      5@     �I@     �s@      N@     Pv@     @g@      v@     �m@      ?@       @     �L@     �W@      @      @     �U@      "@     �e@      L@     @^@     @U@      @       @      A@     �L@      @      @     �J@      @     �^@      <@      V@     �F@                      4@     �B@       @              ?@      @      R@      6@      K@      @@               @      ,@      4@       @      @      6@              I@      @      A@      *@                      7@     �B@                      A@      @      J@      <@     �@@      D@      @              "@      "@                      3@      @      7@       @      .@      7@                      ,@      <@                      .@       @      =@      4@      2@      1@      @      ,@     �d@     �l@      1@      F@      m@     �I@     �f@     @`@     �l@      c@      ;@      �?     �C@      L@      �?      @      I@      @     �U@      <@      T@      D@      @      �?      4@      6@              @      5@      @      I@      .@     �J@      ;@      @              3@      A@      �?       @      =@              B@      *@      ;@      *@              *@     �_@     �e@      0@     �C@     �f@      H@     @X@     �Y@     �b@     @\@      8@      @     �R@     �]@      &@      :@     �a@      6@     �M@     �F@     @W@      N@      (@      @      J@      K@      @      *@      E@      :@      C@     �L@      M@     �J@      (@             �X@     �n@      &@      0@     @]@       @     0�@     �F@     �{@     @Z@      @              O@      e@       @      @     �R@      @      @      <@     �r@      J@      @              N@      e@              @     �Q@       @     �~@      9@     pr@     �I@      @              =@     �Q@              �?      @@       @      c@      3@     �W@      4@       @              ?@     @X@               @     �C@             @u@      @      i@      ?@      �?               @               @              @       @      @      @      @      �?                      B@      S@      "@      *@      E@      @     �b@      1@      b@     �J@      �?              &@       @       @              "@       @     �G@      @      >@      &@                              @       @              @              ;@       @      (@                              &@      @                      @       @      4@      @      2@      &@                      9@      Q@      @      *@     �@@       @     �Y@      &@     �\@      E@      �?              ,@      6@      @      @      *@             �Q@      @     �D@      .@                      &@      G@      @       @      4@       @      @@      @     �R@      ;@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�&�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�i�ĭ=@�	           ��@       	                   �1@�Jф��@�           �@                           @���	��@           �@                           �?+��I@�             r@������������������������       ��'8춆 @�            �o@������������������������       �rI��@             A@                            �?�ko��@�            �s@������������������������       ��sÉ��@t             g@������������������������       �$�G�T�@Q            �`@
                           �?L!���@           ��@                           �?}���Z@�            �r@������������������������       ��Awu@g            �b@������������������������       �\�H��@[            �b@                           @f��"�@C           0@������������������������       �@�I���@9           P~@������������������������       �����@
             ,@                           �?/�%�A@(           ��@                          �<@=��9)@�           `�@                           �?�1nT�b@v           P�@������������������������       �C��H�)@�            �o@������������������������       �wa�@�            �t@                          �>@��O��@;            �X@������������������������       ���W���@#            �I@������������������������       �AO���@            �G@                           @�bv�z�@w           ��@                           �?G;x%Zb	@�           �@������������������������       ��L�~�	@�            �u@������������������������       ��	z
	@�           P�@                           @��gpse@�           ��@������������������������       �zm�$�@;           p@������������������������       ���{�@�            �l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �p@     0�@     �B@     �H@     �|@      T@     �@     @l@     p�@     `v@      =@      @     �P@     `e@      @      "@      _@       @     �~@     @P@     pu@     �\@      @       @      3@     �T@      �?      @     �I@              o@      7@     @a@     �B@                       @      :@              �?      7@             @b@      ,@     �M@      &@                      @      7@              �?      6@             �`@       @     �J@      $@                      @      @                      �?              ,@      @      @      �?               @      &@     �L@      �?       @      <@             �Y@      "@     �S@      :@               @      @      ;@              �?      ,@              O@      @     �G@      7@                      @      >@      �?      �?      ,@              D@      @      @@      @              @      H@      V@       @      @     @R@       @     @n@      E@     �i@     �S@      @              ,@      <@                      ,@      �?     �]@      &@     �U@      ;@                      @      (@                      @      �?      Q@      @      D@      *@                      $@      0@                       @              I@      @     �G@      ,@              @      A@      N@       @      @     �M@      @      _@      ?@     �]@     �I@      @      �?      A@     �L@       @      @     �M@      @     @^@      ?@     �\@     �I@       @       @              @                              �?      @              @               @      *@      i@     �w@      A@      D@     �t@      R@     �}@      d@     ��@     `n@      9@       @     �L@      ]@      @      $@      Q@      @      f@      <@     �d@     �G@      @       @      I@      Y@      @      @     �I@      @     @d@      3@     �c@      =@      @       @      B@      G@      @      @      8@      �?      C@      (@     �P@      2@      @              ,@      K@               @      ;@      @      _@      @     @V@      &@                      @      0@              @      1@      �?      ,@      "@      &@      2@      �?              @      &@               @      @               @              @      0@      �?              @      @               @      *@      �?      @      "@      @       @              &@     �a@     pp@      ?@      >@     �p@     �P@     �r@     �`@      w@     �h@      5@      $@     @V@     �e@      5@      3@      g@      L@      X@      ]@      h@     @]@      0@       @      7@     @P@      &@      @     �N@      4@      ;@      A@     �H@      B@      (@       @     �P@     @[@      $@      ,@     �^@      B@     @Q@     �T@      b@     @T@      @      �?      K@     @V@      $@      &@     �T@      $@      i@      1@     �e@     �S@      @      �?      ?@     �P@      �?       @     �O@      @     �b@      @     �_@      G@      @              7@      7@      "@      "@      4@      @     �I@      $@     �H@     �@@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ&��ThG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���/�N@�	           ��@       	                   �1@�.��@@�           ؠ@                           �?+���N@�           @�@                           �?#�d��@k            �e@������������������������       �W,^��@0            �S@������������������������       ��F�~�4@;            �W@                           @wT,+9j�?&           �{@������������������������       �������?           �z@������������������������       ����Tx%�?	             1@
                            �?ǽ;��%@�           �@                           �?Y��{�@�            �w@������������������������       ���@.Ę @M             `@������������������������       ��}�=@�             o@                            @9��>�@�           ,�@������������������������       ��!h��i@�           ��@������������������������       ����K�@           �{@                           �?��]��@`           t�@                           @'i��Y@�           8�@                          �8@
/���	@            �{@������������������������       �����@y            �f@������������������������       ����@�            pp@                            @px��`�@�            �r@������������������������       �4�H�uo@�             n@������������������������       ���A觑�?%             M@                           @�;�M16	@�           ��@                           �?��NT�
@�           ��@������������������������       ��%;9�@_             b@������������������������       ���@�^
@P           0�@                           @�l�@�             v@������������������������       ��L���@�             k@������������������������       ��Ռ%@N            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     pq@     ��@      >@     �H@     �|@     @X@     Џ@      j@     h�@     0y@      8@      @     �Y@     �s@      &@      0@     @k@      A@     p�@      S@     �~@     �d@      "@      �?      3@      R@      �?      @      K@      @     �q@      .@     �`@      @@              �?      &@      6@      �?              @@      @     �D@       @     �C@      0@                      @      @                      &@      @      8@      @      6@      @              �?       @      0@      �?              5@              1@      @      1@      $@                       @      I@              @      6@             �m@      @      X@      0@                       @      I@              �?      6@             �l@      @      X@      &@                                              @                      "@                      @              @      U@      n@      $@      (@     �d@      ?@     `{@     �N@     v@     �`@      "@              *@     �M@              �?      B@      @      _@      .@      Y@      7@      @              �?      7@              �?       @             �K@      @     �A@      "@                      (@      B@                      A@      @     @Q@      (@     @P@      ,@      @      @     �Q@     �f@      $@      &@      `@      <@     �s@      G@     �o@     @[@      @      �?      I@     �^@      @      @     �O@      2@     �i@      =@     �b@     �Q@      @      @      5@     �M@      @      @     @P@      $@     �[@      1@     @Z@      C@      @      .@      f@     `l@      3@     �@@     �n@     �O@     �r@     �`@     Pr@     �m@      .@      @     �P@     �^@      @      (@     �W@      5@     �`@      F@     �^@     @[@      @      @      E@     �T@      @      @      M@      1@     �G@     �B@     �L@     @T@      @              4@      >@      �?       @      <@      @      <@      @      ?@      9@      @      @      6@      J@      @      @      >@      *@      3@      >@      :@      L@       @      �?      9@     �D@              @      B@      @     �U@      @     �P@      <@              �?      9@     �C@              @      @@      @     �M@      @      H@      6@                               @              �?      @              ;@              2@      @              $@     @[@      Z@      ,@      5@     �b@      E@     �d@     @V@     @e@     @`@       @      $@     @W@     �P@      $@      5@     �Y@     �A@     �R@      R@     @V@     @T@       @              :@      0@              �?      2@              9@      $@      <@      2@       @      $@     �P@     �I@      $@      4@      U@     �A@     �H@      O@     �N@     �O@      @              0@     �B@      @              H@      @     @W@      1@     @T@     �H@                      (@      :@      �?              9@      @     �Q@      $@      H@      5@                      @      &@      @              7@      @      6@      @     �@@      <@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @_�~�c6@�	           ��@       	                   �3@�����@j            �@                           �?�z�6�@�           @�@                            �?..:͂@%           �|@������������������������       ���Hv��@�             o@������������������������       �/a���@�            @j@                           �?������@�            �k@������������������������       �e����� @/             S@������������������������       �h�=�5S@^            @b@
                           �?�Z�{%;	@�           ��@                           �?��5~|@�            �y@������������������������       �\���V�@�            �s@������������������������       ��*��h@<            �X@                            @I�Oj�G	@�           8�@������������������������       ����r�k	@�           `�@������������������������       �o�h7�@            z@                           �?�G-�uq@5           �@                            �?[���r @m           ��@                           �?��A_>@�            �s@������������������������       ���E�M��?v             h@������������������������       ��$�W�@N            �_@                           �?/��?�             p@������������������������       ���h�o�?b            �b@������������������������       ��+>���?G            �Z@                           @���'�@�           �@                            @!���x@           �@������������������������       �bqb��@�           ��@������������������������       ��:����??            �Y@                            �?����@�            �s@������������������������       �OU����@b            �d@������������������������       �qN�F�@a            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �s@     ��@      6@      P@     �z@     @Q@     4�@     �k@     ��@     �t@      ?@      6@     @n@     �u@      *@      G@      t@      K@     �v@     �f@      v@     @l@      <@      @      L@     �X@      @      @      T@      @     �f@     �J@     �^@     �N@      @      @      C@     @R@      @      @     �M@      @     �Y@      D@     �Q@      J@      @      �?      8@     �C@       @      �?      8@      @     �K@      :@     �F@      7@      @      @      ,@      A@       @       @     �A@      @     �G@      ,@      9@      =@      �?              2@      :@               @      5@             @T@      *@      J@      "@                      "@      @                       @              ;@      �?      =@      @                      "@      6@               @      3@              K@      (@      7@      @              1@     @g@     �n@      "@     �D@      n@      H@      f@     @`@      m@     �d@      6@      @      M@      I@       @      $@      C@       @     @V@      5@     @W@      C@      @      @      J@      F@       @      "@      ;@      �?     �F@      1@     @R@     �A@      @              @      @              �?      &@      �?      F@      @      4@      @       @      ,@      `@     `h@      @      ?@     @i@      G@      V@     @[@     `a@     �_@      0@      @     �S@      _@      @      9@     �_@     �@@      K@     �S@     �Q@     �R@      $@      @      I@     �Q@       @      @      S@      *@      A@      ?@     @Q@     �J@      @       @     �Q@      o@      "@      2@     @Z@      .@     (�@     �C@     �z@      Z@      @              &@      V@               @      :@      @     0r@      @     �]@      ;@                      @     �N@              �?      4@      @      c@      @     �K@      2@                      �?      >@              �?      0@             �Y@      @      ?@       @                       @      ?@                      @      @      I@      �?      8@      $@                       @      ;@              �?      @             @a@      @      P@      "@                       @      0@              �?      @             @U@       @      @@       @                      @      &@                      @             �J@      �?      @@      �?               @     �M@      d@      "@      0@     �S@      &@      x@      @@     �s@     @S@      @       @      C@      \@      @      @     �K@      @     �r@      2@     �m@      H@      @       @      B@     @Z@      @      @      E@      @     �p@      2@      h@      G@       @               @      @                      *@              A@             �E@       @      �?              5@      H@      @      &@      8@      @     �T@      ,@      S@      =@                      (@      =@              @      &@       @      B@      &@     �H@      $@                      "@      3@      @      @      *@      @     �G@      @      ;@      3@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�p.hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@����I@�	           ��@       	                   �1@_Bv2�@|           z�@                           @�$�-@{           ��@                           @*"�o-@�            �r@������������������������       ���-=�v@R             `@������������������������       �`��/԰�?k             e@                           @�2L��>@�            �r@������������������������       ���*�@X            ``@������������������������       �������?f            �d@
                           @���s�@           ��@                           �?�6� �l@&           (�@������������������������       �!����@�            �p@������������������������       �d�g�\�@y           ؂@                           �?�����@�           @�@������������������������       ��U@�r@�            �y@������������������������       �4{�w�@�            �v@                           �?��4�@B           0�@                           �?�>����	@           @�@                           �?*6��@�            �k@������������������������       ��e��@/             T@������������������������       �$��Й@c            �a@                          �:@-6�5�+
@�           H�@������������������������       ����O,�	@�            Pw@������������������������       �����	@�            �j@                           @-�{~�@(            �@                           @�WV$@D           8�@������������������������       ��8��@�            `s@������������������������       �pV�И�@             j@                           �?�fj��@�            �u@������������������������       �1�v�Z�@s             f@������������������������       �]�݁�@q            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     @r@     �@      9@      P@      }@     �Q@     D�@     �k@     h�@     0x@     �A@      @      `@     �q@      $@      :@     �o@      C@     X�@     �X@     �~@     �d@      1@              ;@      P@      �?      @     �J@      �?     p@      2@      _@      D@       @              4@      ?@              �?      6@             �a@      @     �H@      7@       @              &@      .@                      2@              F@      @      6@      (@                      "@      0@              �?      @             @X@      �?      ;@      &@       @              @     �@@      �?      @      ?@      �?      ]@      &@     �R@      1@                      @      3@      �?      �?      6@      �?      D@      &@      0@      *@                              ,@              @      "@              S@             �M@      @              @     @Y@     �k@      "@      5@     �h@     �B@     �|@      T@      w@     �_@      .@      @     �N@     @]@      @      ,@     `b@      :@     �d@     �P@      d@     @V@      (@              :@     �B@              �?      8@      @     �Q@      0@      N@      ;@       @      @     �A@      T@      @      *@     �^@      7@     �W@      I@      Y@      O@      $@              D@     �Z@      @      @      J@      &@     `r@      ,@      j@      C@      @              4@     �A@       @      @      E@      @      d@      &@      \@      6@      �?              4@     �Q@      �?      @      $@       @     �`@      @      X@      0@       @      (@     �d@     `l@      .@      C@     �j@      @@     `t@     �^@     r@     �k@      2@      &@     �X@     @]@      $@      =@     @]@      3@     @W@     @R@     �Z@     �]@      .@              5@     �B@              @      A@             �@@      *@      H@      <@       @              ,@      @                      .@              0@              0@      $@       @              @      >@              @      3@              1@      *@      @@      2@              &@     @S@      T@      $@      6@     �T@      3@      N@      N@     �M@     �V@      *@       @     �F@      O@      @      .@     �L@      (@     �F@     �C@     �C@     �D@      (@      "@      @@      2@      @      @      :@      @      .@      5@      4@      I@      �?      �?     �P@     �[@      @      "@     �W@      *@      m@      I@     �f@     @Y@      @      �?      E@      J@      �?      "@      N@      $@     �a@      ?@     @X@      R@      @      �?      &@     �A@              @     �@@       @     @[@      .@      M@     �A@       @              ?@      1@      �?      @      ;@       @      @@      0@     �C@     �B@      �?              8@      M@      @             �A@      @      W@      3@     @U@      =@                      *@      D@                      0@      �?      E@      @      F@      ,@                      &@      2@      @              3@       @      I@      (@     �D@      .@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�mQ;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @=�J��^@�	           ��@                          �2@���XO	@p           
�@                           @�]\�@;           �~@                          �1@�.Y���@4           0~@������������������������       ����A�@�            0p@������������������������       �=��:�T@�             l@������������������������       ���q`�@             &@                           �?�Oo���	@5           \�@	       
                    �?{J�~L)@            �}@������������������������       �����\@�            �l@������������������������       ���{h@�            �n@                           @�@-��
@           ��@������������������������       ����wX�	@�           l�@������������������������       �����	@i            @d@                          �4@w��j��@A           �@                          �1@�LH���@O           ��@                           @늺�s� @�            `x@������������������������       ��K9$l& @�            �s@������������������������       �Q�q'��@-            �S@                            �?�,� K�@`           P�@������������������������       �J��zp�?S            �_@������������������������       �I��*B@           �x@                           @q�\�с@�           ��@                           @���w$@�           ��@������������������������       ����n��@D           ��@������������������������       ���Öj�@�            �p@������������������������       �G�:�L@             5@�t�bh�h5h8K ��h:��R�(KKKK��h��B 
        &@     �r@     �@      B@      K@     �z@     �T@     ȏ@      j@     (�@     �w@      G@      &@      j@     Pt@      =@     �D@     `r@     �N@      x@     �f@     @v@     `o@     �D@       @      8@     �S@       @      @     �P@       @     �a@     �@@      W@     �H@       @       @      8@     �S@       @      @      O@      �?     `a@     �@@     �V@      H@              �?      *@      D@       @      �?      6@             @V@      ,@     �K@      6@              �?      &@      C@               @      D@      �?      I@      3@      B@      :@                                                      @      �?      �?              �?      �?       @      "@      g@     �n@      ;@      C@     `l@     �M@     �n@     `b@     �p@     @i@     �C@             �H@     @R@       @      @     �G@       @     �\@      :@     �V@     �K@      @              4@      ?@       @      @      6@      @     �K@      *@      E@      A@                      =@      E@                      9@      @     �M@      *@      H@      5@      @      "@     �`@     �e@      9@      @@     �f@     �I@     @`@     @^@     �e@     `b@     �A@      @      [@      c@      9@      <@     `c@     �F@      ]@     �W@     `d@     �`@      9@      @      ;@      6@              @      9@      @      ,@      :@      &@      ,@      $@             �W@      k@      @      *@     �`@      6@     ȃ@      =@     |@     �`@      @             �D@     �\@      @      @     �D@      @     py@      (@     `l@     �K@      �?              &@     �F@              @      3@             �f@      @     �Y@      4@      �?              &@      B@              �?      1@             �b@      �?     �U@      $@      �?                      "@              @       @              A@       @      1@      $@                      >@     @Q@      @       @      6@      @      l@      "@      _@     �A@                       @      2@                      @             �Q@      @      5@       @                      6@     �I@      @       @      3@      @      c@      @     �Y@     �@@                     �J@     �Y@      @      @     �V@      2@     @l@      1@     �k@     @S@      @             �E@     �Y@      @      @     @V@      *@      l@      0@     �k@     @S@      @              ;@      R@              �?     �K@      @     @f@      @     @b@     �D@      @              0@      >@      @      @      A@      @     �G@      $@     �R@      B@      �?              $@              �?               @      @      �?      �?      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��TdhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��tV/X@�	           ��@       	                    �?����h�@�           `�@                          �5@é��M�@�           0�@                            �?7y}Ŷ@�            `v@������������������������       ���n��g@F            �\@������������������������       ���P�>@�            `n@                           �?qC��4�@�             r@������������������������       ��$ q�@O            �`@������������������������       ���ƸW�@f            @c@
                           �?�(�O��	@�           ��@                          �4@�m��	@_           @�@������������������������       �Cyc�=@�             l@������������������������       �գm
@�            �v@                           �?A1�0	@�           �@������������������������       �SXTД	@�            �@������������������������       ���MڄZ@�            �o@                           �?T�D	0@'           d�@                          �5@�$�g��@n           8�@                          �3@<q�e @           �y@������������������������       ����Z� @�            0r@������������������������       �]���> @G            �^@                            �?�
+���@l            @e@������������������������       �����5�@            �@@������������������������       ������Q@V             a@                          �7@'���@�           H�@                          �3@\�2H��@�           ��@������������������������       ��5ntI@           �{@������������������������       ��H]=�@�            �w@                           �?�r���5@�             r@������������������������       � ����r@	             .@������������������������       �M.��4�@�            q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     �s@     x�@      :@     �L@     �z@     �R@     �@     �k@     ��@     Pv@     �@@      5@     �k@     pt@      2@     �C@     pr@      M@     �w@     �f@      y@     �o@      >@              R@     �X@      �?      @     @P@      @      c@      7@     �e@      G@      @              4@     �N@      �?       @      >@      @      Z@      &@      Y@      7@      @              @      7@              �?       @       @      =@      @      F@       @                      1@      C@      �?      �?      6@      �?     �R@       @      L@      5@      @              J@      C@               @     �A@              H@      (@     �R@      7@      @              5@      6@              �?      *@              <@       @      >@      &@                      ?@      0@              �?      6@              4@      @     �F@      (@      @      5@     �b@     �l@      1@     �A@     �l@     �K@      l@     �c@     `l@      j@      8@      "@     �C@     �X@      (@      @     �U@      ;@     �R@      N@     �O@      X@      (@       @       @      F@       @             �B@       @     �E@      6@      =@      =@              @      ?@      K@      @      @     �H@      9@      @@      C@      A@     �P@      (@      (@     �[@     @`@      @      <@      b@      <@     �b@     �X@     �d@      \@      (@      (@     �U@     @W@      @      6@     @[@      7@     �W@     @R@     �]@     �V@      (@              8@     �B@              @     �A@      @      K@      :@     �F@      6@              @     @X@      m@       @      2@     ``@      1@     P�@     �C@     @z@     �Y@      @              ;@      S@              @      >@       @     �p@      .@     �`@      :@      �?              0@      H@              @      .@      �?     @l@      &@     �S@      *@      �?              (@      =@                      $@             �c@      "@      O@      &@      �?              @      3@              @      @      �?     @Q@       @      0@       @                      &@      <@                      .@      �?     �E@      @     �K@      *@                              @                      @              &@      �?      @      @                      &@      7@                       @      �?      @@      @      I@      "@              @     �Q@     �c@       @      ,@     @Y@      .@     �u@      8@     �q@     @S@       @              E@      `@      @      $@     �L@      *@     �r@       @      j@     �I@      �?              4@     @P@       @      @      3@             �g@       @     �Z@      ;@                      6@      P@      �?      @      C@      *@      [@             �Y@      8@      �?      @      <@      ;@      @      @      F@       @     �J@      0@     �S@      :@      �?      @      @                                               @       @       @      @                      9@      ;@      @      @      F@       @     �I@      ,@     @S@      7@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@���$�@�	           ��@       	                   �1@&0Y0/<@�           ��@                            �?��L���@�           ��@                           @_{�!R@�            �u@������������������������       �;L��� @�            @o@������������������������       �Y�O,3^@7            �W@                           @�ॢ�@�            �q@������������������������       �[��cp[@`             b@������������������������       ����y��@T            @a@
                           �?y�ǧ@           h�@                           @H�o�@�            �v@������������������������       �1�g�q�@            �i@������������������������       �:��׎>@g            �c@                           �?u���r@&           0~@������������������������       �Wy^	@            �i@������������������������       ���Ƥ�:@�            Pq@                           �?D{�h�@           �@                           �?w�H��	@�           �@                           �?����@           `z@������������������������       ��a˶�@S             _@������������������������       �H��D�l	@�            �r@                           �?�b���	@�            �@������������������������       ���9|@�            `i@������������������������       �B)�I�.
@M           ��@                           @��c���@2           �@                           �?���:;@�             v@������������������������       ��wz��@9            �Y@������������������������       �[�T��@�             o@                           @N0@߻@\            �@������������������������       ����#A�@�           ��@������������������������       �z N�E�@�            �t@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �s@     Ѐ@     �B@      N@      {@     �X@     �@     `o@     X�@     �v@      @@      @     �R@     @f@      @      (@     �`@      1@     �~@     @S@     �u@     �\@      @              7@      T@              �?     �G@       @     �o@      6@     �c@      D@      �?              $@     �I@              �?      2@       @     �a@      &@      V@      6@                       @      >@                      *@             @Y@      @     @T@      *@                       @      5@              �?      @       @      D@      @      @      "@                      *@      =@                      =@              \@      &@     @Q@      2@      �?               @      &@                      *@             @Q@      @      :@      "@      �?              @      2@                      0@             �E@      @     �E@      "@              @      J@     �X@      @      &@      V@      .@     @n@     �K@     @h@     �R@       @       @      0@     �E@       @              F@      @     �]@      ;@      U@      5@               @      (@      9@                      =@      @      F@      9@     �G@      .@                      @      2@       @              .@             �R@       @     �B@      @              @      B@     �K@      @      &@      F@      $@      _@      <@     �[@      K@       @      @      ,@      0@      @       @      =@      @      ;@      8@      D@     �@@       @              6@     �C@       @      @      .@      @     @X@      @     �Q@      5@              (@      n@     �v@      >@      H@     �r@     @T@     �|@     �e@     �|@     �n@      =@      "@     `c@     �f@      6@      ;@      e@      G@     @_@     �[@     �d@     @_@      :@      �?      D@     �N@      @      (@     �P@      .@     �R@      ;@     @Q@     �F@       @      �?      0@      (@                      ;@              =@       @      ?@      @       @              8@     �H@      @      (@      D@      .@     �F@      9@      C@     �D@      @       @     �\@      ^@      3@      .@     @Y@      ?@     �I@     �T@     �W@      T@      2@             �A@     �F@      @      @      7@              0@      4@      <@      6@      @       @      T@     �R@      ,@      "@     �S@      ?@     �A@     �O@     �P@      M@      .@      @     @U@     `f@       @      5@     ``@     �A@     u@      P@     �r@     �^@      @              7@     �J@      @      "@     �C@      0@     �R@      =@      P@      D@      �?              @      (@              �?      ,@      @      F@       @      4@       @                      2@     �D@      @       @      9@      *@      >@      ;@      F@      C@      �?      @      O@     �_@      @      (@      W@      3@     pp@     �A@      m@     �T@       @      @     �A@      R@      �?      @      K@      @     �g@      6@      e@      H@      �?              ;@      K@      @      "@      C@      (@     @R@      *@      P@      A@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�_t1f@�	           ��@       	                    �?�.�ӫR@           ��@                          �5@�H��f�@A           �@                            �?LS�q�@�            �p@������������������������       �B<9Z��@-            @U@������������������������       �ֶ���@t            �f@                           �?�SаB�@�            `n@������������������������       �Ē[�g@8             U@������������������������       �wnL�E@h            �c@
                            �?��Uo��@�           8�@                           @���� �?t            `h@������������������������       ��	�#�8�?J            @_@������������������������       �ߕi�?*            �Q@                           @Om^\4@V            �@������������������������       ��-�_�@N             ^@������������������������       �n��?@           �z@                          �3@Ψ^�f@�           Ȥ@                           @~Vݛ�@:           X�@                           @�=�O�@e            �c@������������������������       �i�U{��@:            �V@������������������������       ���+�@+            �P@                           �?�]���@�           p�@������������������������       �|��U�@�            �k@������������������������       �,� ���@@           @                          �9@?s��	@j           �@                            �?K�7��c@           ��@������������������������       ���P�g@�            �s@������������������������       ��q<@6           x�@                           @�v����	@e           x�@������������������������       �{��c
	@V             a@������������������������       ��ir�Or	@           p|@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@      t@     Ȁ@      A@      J@      }@     @V@     ��@     �j@     h�@     @v@      ?@      �?     @W@     �c@      @      @     �[@      @      }@      H@     �q@     �Q@      @      �?      J@     �S@      @      @     @P@      @     �Z@     �@@     �]@      E@      @              .@      C@              �?      :@      @     �S@      1@      R@      .@      �?               @      1@                      @              <@      @      :@      �?                      *@      5@              �?      6@      @     �I@      $@      G@      ,@      �?      �?     �B@      D@      @      @     �C@              ;@      0@     �G@      ;@      @      �?      ,@      $@                      0@              3@       @      .@      @       @              7@      >@      @      @      7@               @      ,@      @@      6@      �?             �D@     �S@      �?       @      G@      @     `v@      .@      e@      =@      �?               @      ,@      �?              0@      �?     �[@       @     �C@       @      �?               @      "@                      @      �?      P@              A@      @      �?                      @      �?              "@             �G@       @      @      �?                     �C@      P@               @      >@      @     �n@      *@      `@      5@                      2@      @                      (@      �?     �H@      @      4@       @                      5@     �M@               @      2@       @     �h@      @     @[@      *@              1@     �l@     �w@      >@      G@     v@     �T@     8�@     �d@     �~@     �q@      :@      @     �E@     �_@      @       @     �T@       @     @q@      H@     �f@     �U@      @      @      $@       @               @      5@      �?     �G@      3@      @@      ,@              @      @      @              �?      0@              ,@      .@      2@      *@                      @      @              �?      @      �?     �@@      @      ,@      �?              �?     �@@     �]@      @      @     �N@      @     �l@      =@     �b@      R@      @      �?      4@      :@      @      @      >@      @     �E@      1@      ?@     �A@      @              *@      W@      @       @      ?@      �?     @g@      (@      ^@     �B@              *@     @g@     �o@      8@      C@     �p@     �R@     0q@     �]@     ps@     �h@      5@      @      ]@     �h@      *@      =@     �f@     �@@     �j@      L@     �k@     @\@      (@              G@     �H@      @      "@      F@      @     �M@      3@     �G@      <@      @      @     �Q@     �b@      $@      4@     @a@      ;@      c@     �B@     �e@     @U@      @      @     �Q@      L@      &@      "@     @V@     �D@     �O@      O@     @V@     �U@      "@      �?      1@      .@      @              &@      (@      @      ;@      5@      3@      @      @     �J@     �D@       @      "@     �S@      =@     �M@     �A@      Q@     �P@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���xhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�����x@�	           ��@       	                     @U!1vth@
           H�@                           �?�&�և@<           X�@                            �?u�ػ?4@           �{@������������������������       ���%�x�@�            �t@������������������������       ���%�@I            @]@                            �?S>�x�8@           �|@������������������������       ����g�@s            �g@������������������������       �^�6͸[@�            �p@
                           �?����@�            pt@                           �?�m��@s            �f@������������������������       ���x���@;            @V@������������������������       �)�n29@8            �W@                           @k)k5 �?[             b@������������������������       ����I.\ @*            �N@������������������������       ���P��?1            �T@                           @��?��p@�           �@                          �4@�b��	@�           \�@                           �? ���?@w           ��@������������������������       �z�ۥ&�@t            @g@������������������������       �,�+s��@           @z@                            @<�("n�	@f           ȍ@������������������������       �Dz*k�	@z           ��@������������������������       �����,�	@�            Pv@                           @uKsi2k@�           ��@                           @:.4��@�           �@������������������������       �Ԋbm��@�           p�@������������������������       ��Sğ@�            @s@                            �?_���I@             >@������������������������       ���	M�1@	             0@������������������������       �RM棿@
             ,@�t�b�N      h�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     ȁ@     �B@     �P@     �|@     @T@     ��@      k@     H�@     �u@     �C@      �?     �T@     �d@      @      @     @\@      "@      |@     �C@     �q@     @Q@      "@      �?      K@     @]@      @      @     �U@      "@     @t@      7@     �k@      L@      "@      �?      6@      M@       @       @     �H@      @     �g@      ,@     @Q@      >@      @      �?      2@     �D@       @       @      E@      @     �`@      $@     �F@      <@      @              @      1@                      @      @      L@      @      8@       @                      @@     �M@       @       @     �B@      @     �`@      "@     �b@      :@      @              "@      A@       @              1@       @      H@      @      N@       @      @              7@      9@               @      4@      �?     @U@      @     �V@      2@       @              =@     �G@               @      ;@             �_@      0@     �P@      *@                      4@     �E@               @      2@             �F@      .@      =@      &@                      "@      2@              �?      &@              6@      @      .@      @                      &@      9@              �?      @              7@       @      ,@      @                      "@      @                      "@             @T@      �?      C@       @                      @      @                      @              >@      �?      .@      �?                      @                              @             �I@              7@      �?              (@     @k@     Py@     �@@      N@     �u@      R@     ��@      f@     P�@     Pq@      >@      (@     @b@     �m@      7@      G@     @o@     �K@     �h@     @b@     �l@     �g@      ;@       @     �A@     �U@      @      $@     �W@      "@     �Z@      M@     �[@     @S@      (@       @      &@      <@      @              ?@      @     �B@      9@      4@      7@                      8@      M@      �?      $@     �O@      @     �Q@     �@@     �V@      K@      (@      $@     �[@      c@      2@      B@     �c@      G@     �V@      V@     �]@      \@      .@      @     �P@      U@      @      @@     @Z@      @@     �F@      L@     �S@     �S@      @      @     �F@      Q@      (@      @     �I@      ,@      G@      @@      D@      A@       @              R@     �d@      $@      ,@     �W@      1@     �t@      ?@     Pr@      V@      @             �P@     �d@      $@      $@     �V@      *@     �t@      <@     �q@      V@      @              J@     �]@              @     �Q@      @     q@      5@     @h@     �E@       @              .@     �G@      $@      @      4@       @      L@      @      W@     �F@      �?              @      �?              @      @      @      �?      @      @                              �?                      @      �?      @              �?      @                              @      �?                      @              �?       @       @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJE�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�ct�[U@�	           ��@       	                    �?�y���@m           6�@                           �?�S��g@�            �@                           �?H2�ç.@1           `~@������������������������       �r���5�@m            @f@������������������������       ��˜�@�            @s@                            �?1�≩�@m            @g@������������������������       ��Ǳ @$            �Q@������������������������       ��B�@I            �\@
                           �?���Zt	@�           �@                           �?��d!)�	@�           H�@������������������������       ��
g?@           �{@������������������������       ��Jr�"
@�           ��@                          �5@�=��'o@           �z@������������������������       ��1W&[p@�            �k@������������������������       �(�8m�q@�            `i@                          �5@��<J�>@K           ��@                          �4@s��s3�@�           �@                           @�s|�@X            �@������������������������       �w��1H@�            �j@������������������������       �M�(XT�@�           h�@                           @%��@��@i            �c@������������������������       ��yfp@J            �[@������������������������       �c��H�@             H@                          �7@.E�p2@�           `�@                           @����@�            �m@������������������������       ����6�@<            �Z@������������������������       �tr��<�@Q            @`@                           @� ��>@�             x@������������������������       �s�$I@�             k@������������������������       ���z�;�@g            �d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      r@     ��@      :@     �P@      }@      R@     ��@     �j@     X�@     �w@     �@@      .@     @j@      t@      4@     �I@     �s@      K@     �w@     `e@     �w@     p@      >@             �P@     @W@       @      $@     �T@      @     �e@     �@@     @b@      M@      @              L@     �S@       @       @     @P@      @     �X@      >@     �W@     �H@      @              9@      7@                      6@             �J@       @      E@      &@                      ?@     �K@       @       @     �E@      @     �F@      <@      J@      C@      @              &@      .@               @      1@             �R@      @      J@      "@       @              �?      @               @      @              <@              :@      �?       @              $@       @                      *@             �G@      @      :@       @              .@     �a@     `l@      2@     �D@     `m@     �I@     `i@     @a@     �m@     �h@      9@      .@     �[@     �c@      *@      =@     `f@      C@     �^@     �W@     �d@     �c@      7@             �B@     @P@      �?      0@     �Q@       @      R@      =@      T@      L@      @      .@     @R@     �W@      (@      *@      [@      >@      I@     �P@     �U@     @Y@      0@             �@@      Q@      @      (@      L@      *@     @T@     �E@     �Q@      E@       @              "@     �B@      @       @      7@      @      M@      4@     �C@      2@                      8@      ?@              @     �@@       @      7@      7@      ?@      8@       @      �?      T@      n@      @      0@     �b@      2@     Ȃ@     �D@     �z@     @_@      @             �B@     `c@      �?      *@     �O@      $@     �|@      1@     0q@     �M@       @              B@      `@      �?      "@      F@      @     Py@      .@     �m@      J@       @              .@      D@                      "@      @     �R@      @     �J@      2@                      5@      V@      �?      "@     �A@      �?     �t@      (@     �f@      A@       @              �?      ;@              @      3@      @     �J@       @     �C@      @                      �?      2@                      &@      @     �C@      �?      ?@      @                              "@              @       @      �?      ,@      �?       @      @              �?     �E@     �U@      @      @     �U@       @     �a@      8@     @c@     �P@      �?              .@     �K@      @      �?      ;@       @     �L@       @      I@      8@                      "@      ;@                      @      �?      C@      �?      3@       @                      @      <@      @      �?      8@      �?      3@      �?      ?@      0@              �?      <@      ?@       @       @     �M@      @     �U@      6@      Z@      E@      �?      �?      ,@      7@              �?      C@              J@      $@      M@      3@      �?              ,@       @       @      �?      5@      @      A@      (@      G@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJC�-'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�����6@�	           ��@       	                    �?����@b           0�@                           �?BR�(gt@�           ��@                          �4@NZu� 2@�            �r@������������������������       �O�S�05@�            `m@������������������������       �D=���]@$            �P@                           �?���9@.            }@������������������������       �b�W�P}@V            �`@������������������������       ���kX�@�            �t@
                           @�%l[�@�           h�@                          �3@�bm�@�             u@������������������������       ��'~eQ@�             n@������������������������       ��>�p��@D            @X@                           @s���_�@�            �@������������������������       �K	 �ѝ@�            �q@������������������������       �����:v@           ��@                           @8A�<Y[@=           Ě@                           �?l^�p% 	@�           4�@                           �?� �WI	@           ��@������������������������       ����B�@�             r@������������������������       ���i�xm	@e           �@                          �=@_h�Q�@�            �m@������������������������       ���A9f+@�             j@������������������������       �2j`	�@             >@                          �7@_��}�@�            �@                           @�
s2[�@�            �k@������������������������       ��G��w@_             c@������������������������       �2�ha9�@/             Q@                           �?�G�ޫr@�            �x@������������������������       �x��&w�@J             _@������������������������       �#gT�@�            �p@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     @t@     0�@      A@     �H@     p|@      N@     �@     �k@     ��@      v@      @@      "@      a@     �s@      *@      :@     @k@      8@     H�@     �Y@     �|@     �c@      0@      "@      M@     �\@      @      2@      ^@      $@     �b@      P@     �_@     @T@       @      @      3@      K@      @      @      K@      @      N@      >@     �A@      >@      �?      @      "@      B@      @       @     �F@      �?      K@      ;@      :@      <@      �?      �?      $@      2@      @      @      "@       @      @      @      "@       @              @     �C@      N@              *@     �P@      @     �V@      A@     �V@     �I@      @              &@      5@                      &@              D@      @      =@      0@              @      <@     �C@              *@     �K@      @     �I@      =@      O@     �A@      @             �S@     �i@      @       @     �X@      ,@     ��@     �C@     u@     �S@       @              7@      G@      @      @      >@      @     �Y@      3@     �S@      >@                      5@      A@              �?      ,@             �R@      *@     �O@      5@                       @      (@      @       @      0@      @      <@      @      0@      "@                      L@     �c@      @      @      Q@      &@     �|@      4@      p@      H@       @              6@     �J@                      *@      "@     @Z@      @     �N@      "@      @              A@     �Z@      @      @     �K@       @     0v@      0@     �h@     �C@      @       @     `g@     pp@      5@      7@     �m@      B@     �s@     �]@     Pr@      h@      0@      @     �b@      f@      3@      3@     �e@      ;@     �a@     �W@     �b@     �`@      0@      @     @^@      a@      3@      1@     @b@      4@     �W@     �Q@     �[@     @[@      ,@      @     �A@      G@       @      @     �I@      @     �F@      7@     �C@     �@@      @      @     �U@     �V@      1@      ,@     �W@      0@     �H@     �G@     �Q@      S@      "@              ;@      D@               @      ;@      @      G@      9@     �C@      7@       @              7@     �B@               @      7@      @      E@      2@      B@      7@      �?              @      @                      @      @      @      @      @              �?      �?     �C@     �U@       @      @      P@      "@      f@      8@      b@     �N@                      3@      F@       @              4@      @     @Q@      @     �B@      7@                      1@      <@      �?              &@      �?     �L@      @      5@      *@                       @      0@      �?              "@       @      (@              0@      $@              �?      4@     �E@              @      F@      @      [@      5@     �Z@      C@                      �?      1@                      "@      @     �D@      @     �C@      "@              �?      3@      :@              @     �A@      �?     �P@      2@      Q@      =@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�B�mhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?/?{6<@�	           ��@       	                   �<@|KNn@�           ��@                            �?����i�@�           p�@                          �8@G5�~��@�            �r@������������������������       �9�|}$�@�             o@������������������������       ���~���@              J@                          �3@���ԛ�@           x�@������������������������       ��ە�u@�            �w@������������������������       �n4��@           @{@
                           @'at�c�@@            �X@                          �=@���R�[@-            �Q@������������������������       ���aU��?             >@������������������������       �%��N�@            �D@                           @������ @             <@������������������������       �� �P��?	             *@������������������������       ���\�O� @
             .@                           @bw�� @�           �@                           �?)2{�b	@�           ܗ@                           �?�
ƨ/�	@�           ��@������������������������       �OP[���@           �y@������������������������       ��?�G�
@�           h�@                           �?;OX�	*@           y@������������������������       �g��Azj@            �@@������������������������       ��Z��@�             w@                          �7@��0�@�           L�@                           @O�3���@           ؊@������������������������       ���ҹ�-@�           H�@������������������������       ��8N�'@�            @j@                           @�Lb��4@�            �s@������������������������       �3J���@t             g@������������������������       �إE���@N            �_@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     �@      =@     �H@      |@     �S@     ��@      n@     ��@     �t@      @@      �?     �T@     �c@      @      @     @X@      @     0{@     �F@     �q@      W@      @      �?      S@     �a@      @       @     �U@      @     `z@     �C@      q@      P@      @      �?      0@      =@                      9@      @     @\@      @     �V@      1@      �?              (@      8@                      8@       @     �Z@      @      Q@       @      �?      �?      @      @                      �?      �?      @       @      6@      "@                      N@     @\@      @       @     �N@       @     Ps@     �@@     �f@     �G@      @              .@      @@                      <@       @     �d@      .@     @W@      <@      �?             �F@     @T@      @       @     �@@              b@      2@     @V@      3@       @              @      ,@              @      &@              *@      @      ,@      <@       @              @       @              @      "@              @      @      @      9@       @              �?      @                       @                              @      3@                      @      @              @      @              @      @      @      @       @                      @                       @              $@              @      @                               @                                      "@              �?      �?                              @                       @              �?              @       @              *@      k@     pz@      :@     �E@     v@     �R@     �@     �h@      �@     @n@      :@      (@     �c@     @l@      5@      B@     `n@      M@      h@     `b@     �n@      e@      4@      (@      _@     �b@      4@      9@     `g@      F@      ]@      ]@      g@     �`@      0@       @      @@      O@      �?      "@     @P@      &@     �K@      B@     �V@     �F@      �?      $@      W@      V@      3@      0@     �^@     �@@     �N@      T@     �W@     �U@      .@              A@      S@      �?      &@      L@      ,@     @S@      ?@     �N@      B@      @               @      @               @      @      �?       @      @       @      @                      @@     �Q@      �?      @     �J@      *@     �R@      :@     �M@      @@      @      �?     �M@     �h@      @      @     �[@      0@     �w@     �H@     �p@     �R@      @             �B@     �c@      @      @      O@      *@     �r@      1@     `j@      H@      @              =@      \@      �?      �?     �D@      @      n@      *@     �d@     �C@      @               @     �G@       @       @      5@       @     �N@      @     �G@      "@      �?      �?      6@      C@       @      @      H@      @     �S@      @@      L@      :@       @      �?      "@      7@               @     �B@              M@      &@      =@      *@       @              *@      .@       @       @      &@      @      4@      5@      ;@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�P�ɹy@�	           ��@       	                    @�#>+�,@�           ʥ@                           �?U1����@k           ,�@                           �?���X�@           �y@������������������������       �<����@�             i@������������������������       �E-c?v@�            �j@                          �4@ED�K	@[           `�@������������������������       �f�ٯut@�            �v@������������������������       �bC<N�	@s            �@
                          �4@K���Ew@�           h�@                          �0@����s@�           x�@������������������������       �x���{&�?A            @Y@������������������������       �c���@�           P�@                           �?c.���@�           X�@������������������������       ���6*�@�            �t@������������������������       �]4l8��@�            �s@                           �?L�?>�@�           ��@                           �?8�7j�@�            `u@                           �?v2�ū�@~             i@������������������������       �*�#�*@C            @Z@������������������������       �'"�2��@;            �W@                           @�ِ�a��?T            �a@������������������������       ��-��> @            �E@������������������������       �Bh�g�h�?;            �X@                           �?K����@�           p�@                           �?0^w�m@(             P@������������������������       �3�t��H@             3@������������������������       ������@            �F@                           @6�ߔo�@�           p�@������������������������       ��P��/�@�            �s@������������������������       ��o~��R	@�            y@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     r@     x�@      =@     �K@     P~@     �W@      �@     �j@     h�@     `x@     �A@      "@      g@     �w@      .@     �C@     �t@     @P@     ��@      d@     ��@     pp@      :@      "@     @\@     �e@      $@      5@     �i@     �G@      l@      _@     `m@      e@      6@       @      B@     �L@      �?      @      L@      @     �Y@      ,@      Y@      ?@      "@       @      1@      ;@      �?      @      <@      @      J@      &@      @@      6@      �?              3@      >@                      <@              I@      @      Q@      "@       @      @     @S@     �]@      "@      2@     �b@     �E@     �^@     �[@     �`@      a@      *@              4@     �F@      @              L@      @      S@     �F@     �I@      J@      @      @     �L@     @R@      @      2@     �W@      C@      G@     @P@      U@     @U@      @             �Q@     �i@      @      2@     �_@      2@     @      B@     pv@     �W@      @              ?@     @Y@      �?      $@      G@      @     �u@      0@     @f@     �E@      �?              �?      6@                      @              G@              7@      @                      >@     �S@      �?      $@     �D@      @     s@      0@     `c@     �C@      �?              D@     �Y@      @       @     @T@      *@     @b@      4@     �f@      J@      @              6@     �L@      �?      @      G@       @     �P@      @     �W@      7@      @              2@      G@      @       @     �A@      @      T@      .@     �U@      =@               @     @Z@     �b@      ,@      0@     �b@      >@     `n@      K@     `k@     �_@      "@              ;@      D@       @      @      D@       @      ^@      *@      Q@      :@                      7@      C@       @       @      <@       @      E@      &@     �A@      1@                      "@      (@       @      �?      3@       @      4@      "@      8@      @                      ,@      :@              �?      "@              6@       @      &@      $@                      @       @               @      (@             �S@       @     �@@      "@                                                      @              3@       @      @       @                      @       @               @      @             �M@              :@      �?               @     �S@      [@      (@      (@     �[@      <@     �^@     �D@     �b@     @Y@      "@              @      &@                      *@       @              .@      @       @       @                      "@                      �?      �?               @      �?      @       @              @       @                      (@      �?              *@      @      @               @      R@     @X@      (@      (@     �X@      :@     �^@      :@      b@     @W@      @      @      8@     �H@      @      �?      H@      @      Q@       @     @P@     �D@      �?       @      H@      H@      @      &@      I@      4@     �K@      8@     �S@      J@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�2-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              �?��~L�J@�	           ��@       	                    �?*��b@7           ~�@                           @+K���@�           ��@                          �;@�
�k�@�            �w@������������������������       �՚��}@�            0u@������������������������       ��Q��^@            �D@                           @T�.�t�@�            0t@������������������������       �8�һ� @b            �e@������������������������       ���9<@e            �b@
                           @np��0@�            �@                          �5@�`1�)n	@�           Ј@������������������������       ���< �4@�            �x@������������������������       �7pݑ��	@           y@                           @�G�lm@�           0�@������������������������       �X��4�@�            v@������������������������       �n�}�g@�            Pp@                          �5@�S� @a           (�@                          �1@L���B|@\           ��@                          �0@m��0_@�            �p@������������������������       �B��$B&@*            �N@������������������������       ��6%�S@�            �i@                           �?���(� @�           `�@������������������������       ���1��@�            `m@������������������������       ��Q�a*�@            ~@                            @�9,
O@           ��@                           @�A���4@�             q@������������������������       �m�8�C�@s            �g@������������������������       ����J�@7            �T@                           �?a�+�a�@[           �@������������������������       �x����>	@�            �u@������������������������       �\���v@|            �h@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �r@     �@     �@@     �J@     p~@     �T@     ؎@     `k@     ��@     �u@      5@      @     �e@     �r@      0@      @@     �m@      G@     �@     @]@     �{@     �i@      ,@       @     �K@      \@       @      @      P@      �?     �l@      7@      c@      J@      @       @     �F@      G@      �?      @      G@      �?     @W@      2@     @U@      A@      @             �D@     �C@      �?       @      G@              W@      *@      T@      6@      @       @      @      @               @              �?      �?      @      @      (@       @              $@     �P@      �?              2@             @a@      @     �P@      2@                       @      D@                      �?             @S@      @      @@      &@                       @      :@      �?              1@             �N@             �A@      @              @      ^@     �g@      ,@      <@     �e@     �F@     �q@     �W@     pr@      c@      "@      @     �T@     @]@      &@      5@      ]@      B@     @W@     @R@     �_@     @Z@       @             �B@      Q@      @      @      E@      ,@     �N@      ;@     @R@      M@       @      @      G@     �H@      @      ,@     �R@      6@      @@      G@     �J@     �G@      @             �B@     @R@      @      @     �M@      "@     `g@      5@      e@      H@      �?              (@     �E@      @       @      D@      @     �Z@      $@      Z@      9@                      9@      >@              @      3@       @      T@      &@     @P@      7@      �?      (@     @_@     Pq@      1@      5@      o@      B@     �}@     �Y@     Pu@     �a@      @      @      G@     `c@      @      @     �[@      0@     `u@     �H@     �f@      O@      @              .@     �D@      @              4@             @\@      *@     �I@      $@       @              @      $@                      @              9@              &@      @                      (@      ?@      @              *@              V@      *@      D@      @       @      @      ?@     �\@      @      @     �V@      0@     �l@      B@     �`@      J@      @              ,@      ;@               @      1@       @     �Y@      @      J@      (@              @      1@     �U@      @      @     @R@      ,@     �_@      >@      T@      D@      @      @     �S@     �^@      &@      0@     @a@      4@     �`@     �J@     �c@     �S@       @      @      7@      D@      �?      @      N@      @      H@      *@     �K@      1@              @      2@      9@      �?      @      >@      @     �B@      @     �F@      (@                      @      .@                      >@              &@      @      $@      @              @      L@     �T@      $@      $@     �S@      ,@     �U@      D@     �Y@     �N@       @      @      F@      N@      "@       @      K@      (@      :@     �@@      N@      C@       @              (@      6@      �?       @      8@       @      N@      @     �E@      7@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�F41hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?��2�`@�	           ��@       	                   �<@�}ͫK�@�           D�@                           �?������@�           ��@                           �?��e��@�            `x@������������������������       �ꢄj�@b            �a@������������������������       �OOƐ�@�            �n@                           @���*@�           �@������������������������       �pV�?�@�            �q@������������������������       ���6�	�?�            �x@
                            �?%����@>            @Z@������������������������       �5��܁�@             ;@                           @�U!g�3@.            �S@������������������������       ��^�/@#             N@������������������������       �Rq��mZ�?             2@                            @�m=�V;@�           p�@                           @��Q�@�           0�@                          �3@�����U	@Z           ��@������������������������       ���X��@�            �p@������������������������       �ǵ[���	@�           H�@                          �<@ɪe�i�@k           Ѝ@������������������������       ��w��	�@K           H�@������������������������       �
 aC@             �H@                           �?b�V�}	@�           `�@                          �8@z��|s	@5             U@������������������������       �U�mp�d@             F@������������������������       ����9@             D@                           @�r���@�           ��@������������������������       �y�E��@           �|@������������������������       �='�E�	@�             q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        7@     q@     @�@      >@      J@      }@      U@     �@      p@     @�@     @u@      B@       @     �P@     �b@      @      &@     �[@      $@     0{@      F@     0p@     @R@      @       @     �M@      a@      @       @     �W@       @     @z@     �A@     �n@      H@       @       @      A@     �O@      @      @     �G@      @      Y@      =@      S@      =@      �?       @       @      ,@                      &@             �M@      @      A@      $@                      :@     �H@      @      @      B@      @     �D@      8@      E@      3@      �?              9@     @R@      �?      @      H@      @      t@      @     `e@      3@      �?              1@      A@              @      =@      @     @Z@             @T@       @                       @     �C@      �?       @      3@             �j@      @     �V@      &@      �?               @      (@              @      0@       @      .@      "@      (@      9@      @               @      @                       @       @      �?      �?      @       @      @              @      @              @       @              ,@       @      "@      7@                      @      @              @       @              @       @      @      6@                              @                                      @              @      �?              5@     �i@     @w@      :@     �D@     v@     �R@     p�@     �j@     (�@     �p@      ?@      &@     �b@      p@      (@      9@     `o@     �J@     �{@     �a@     �x@     `e@      2@      &@     @V@     @_@      @      3@     `d@     �E@     �b@     �Z@      b@     �Z@      .@      �?      0@      <@      �?             �A@      @      S@      B@      E@      5@      @      $@     @R@     @X@      @      3@      `@     �B@      R@     �Q@     �Y@     �U@      (@              O@     ``@      @      @      V@      $@     �r@     �B@      o@      P@      @             �G@     �^@      @      @     �S@      $@     �r@     �A@     �n@     �L@      @              .@       @      �?              "@               @       @      @      @              $@     �K@      ]@      ,@      0@     �Y@      5@     �a@     �Q@     `c@      X@      *@       @      @      ,@              @      &@      @       @      0@      *@      $@      @      �?       @      $@              @      &@      �?              @      @      @              �?      @      @                               @       @      $@      @      @      @       @      I@     �Y@      ,@      *@     �V@      2@     �a@     �K@     �a@     �U@       @      @      >@      L@      @      @     �K@      "@      W@      8@     @[@      N@      @      @      4@      G@      @       @      B@      "@     �H@      ?@     �@@      :@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���KhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @D��74N@�	           ��@       	                    �?�7�$�@u           `�@                            �?/�����@           (�@                           �?Sq�)��@�             o@������������������������       ��KkVXD@1            �T@������������������������       ����<�@d            �d@                            @fS�9��@y           `�@������������������������       ����Φ)@�            0p@������������������������       �jq�"��@�            �t@
                           �?��ϳh�@g           ��@                          �<@��î�@�            0v@������������������������       �]�s2�@�            �s@������������������������       �޸��`�@            �B@                          �<@�6��x	@�            �@������������������������       �����u	@?           P�@������������������������       ������@I            �_@                           �?t:��@!           d�@                           @�W"�� @]           x�@                          �4@2�=^Sz�?�            �v@������������������������       ��xR�*6�?�            0p@������������������������       � �0�b@E            �Z@                            @/�&�q_@z            @h@������������������������       �
��^�@[            �b@������������������������       �l(Ʋ��?            �F@                          �7@KG��Q�@�           ��@                           @v\ 9@	           ��@������������������������       �����M>@�            �@������������������������       ��:'i`(@�            �j@                            �?&z�	��@�             s@������������������������       ���o�@_            �c@������������������������       ��|r)ˢ@\            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@     �r@     ��@      4@      K@     �{@     �T@     8�@     �i@      �@     �w@      B@      6@     �i@      v@      0@     �D@     �r@     @Q@     w@     �e@     �w@     �p@      >@      &@     �R@      b@      (@      @     �[@      ;@      c@     �O@      _@     @Z@      @              (@      F@               @     �@@      @     �P@      7@     �B@      5@      @              @      ,@                      2@      @      7@      @      *@      �?      �?              "@      >@               @      .@       @     �E@      2@      8@      4@      @      &@     �O@      Y@      (@      @     �S@      4@     �U@      D@     �U@      U@      @      �?      >@      G@      �?      �?      >@      &@      >@      =@      B@     �E@      �?      $@     �@@      K@      &@      @      H@      "@      L@      &@     �I@     �D@       @      &@     �`@      j@      @     �A@      h@      E@      k@     �[@     �o@      d@      7@              A@      N@                      C@      �?     �S@      1@      V@      A@      @             �@@      K@                      B@      �?     �R@      *@      U@      4@       @              �?      @                       @              @      @      @      ,@      @      &@     �X@     �b@      @     �A@     @c@     �D@     `a@     �W@     �d@     �_@      2@      &@     @U@      a@      @      ?@      a@      B@     �`@     �S@      b@     �W@      0@              *@      (@              @      1@      @      @      0@      4@      @@       @      �?      W@      k@      @      *@     �a@      *@     ��@      @@     �z@     �]@      @              ,@     �Q@      �?              8@      @     �p@      @     @a@      >@                      "@      F@                      .@      @     �h@             �T@      ,@                       @      =@                      @             `c@              M@      @                      �?      .@                      $@      @      E@              8@      $@                      @      ;@      �?              "@      �?     �R@      @      L@      0@                      �?      :@      �?               @      �?     �G@      @     �F@      0@                      @      �?                      �?              ;@      �?      &@                      �?     �S@      b@      @      *@      ]@       @     pv@      ;@     �q@      V@      @             �E@     �^@              &@     �Q@      @      r@      1@     @i@      M@      @              A@      X@               @      F@      @     �l@      (@      c@      C@       @              "@      ;@              "@      ;@      @     �M@      @      I@      4@       @      �?     �A@      6@      @       @     �F@      �?     �Q@      $@      U@      >@       @              ;@      0@                      ,@      �?     �@@      @      G@      ,@              �?       @      @      @       @      ?@              C@      @      C@      0@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ==hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��XXxf@�	           ��@       	                   �8@����@u           >�@                           �?���@�           8�@                           �?��EA0@!           P|@������������������������       ��[
�@�            �t@������������������������       ����B�@U             _@                            @�Z>�@�           $�@������������������������       ���%9�@�           ؄@������������������������       ��X4�K@@           �z@
                           @��D��	@�           ��@                           �?��9j�	@o           0�@������������������������       ���_�Ƶ@Z            @b@������������������������       ��?*�L�	@           @{@                          �:@�Zej#@+            �R@������������������������       �D
$[�@             8@������������������������       �N	�y"@            �I@                            �?�l�,@@           ��@                           @��F�@�            �x@                          �7@�<�@�            �m@������������������������       �YŌ)�+�?�            �h@������������������������       ��[OS@             C@                           �?Y6Jj��@]            `c@������������������������       ���z �_@-             S@������������������������       ��4X�	P @0            �S@                          �7@��&˼�@F           ��@                           @0J3�ԉ@�           �@������������������������       �鄿�W�@�             m@������������������������       �����}�@�           ��@                           @?y߸3P@�            t@������������������������       ��guFi@Y            �a@������������������������       �����@e            @f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     s@     p�@     �A@     @P@     �{@      S@     x�@     �j@     (�@     �u@      ?@      5@     @k@     �t@      5@      H@     �s@      M@      x@      g@     �w@     �k@      ;@      *@     �`@      l@      *@      ;@     �m@      @@     pt@     @Y@     �r@      `@      0@             �E@     �K@      �?      @      J@      @     �a@      3@     @Z@      ;@       @              >@      I@      �?       @      F@      @     @T@      2@      T@      2@       @              *@      @              �?       @              O@      �?      9@      "@              *@     �V@     @e@      (@      8@      g@      =@      g@     �T@      h@     @Y@      ,@      @      P@     @X@      @      ,@      W@      6@      ]@     �N@     �^@      M@      &@      @      ;@     @R@       @      $@     @W@      @      Q@      5@     �Q@     �E@      @       @      U@     �Z@       @      5@     �S@      :@     �L@      U@     �T@      W@      &@      @     @R@     @X@       @      5@      R@      7@     �I@      O@      T@      T@       @      @      ,@      :@               @      7@      @      5@      &@      5@      2@      �?       @     �M@     �Q@       @      3@     �H@      3@      >@     �I@     �M@      O@      @      �?      &@      "@                      @      @      @      6@       @      (@      @              @      @                               @       @      @       @      �?       @      �?      @      @                      @      �?      @      1@              &@      �?      �?     �U@     `l@      ,@      1@     �`@      2@     x�@      =@     �z@      `@      @              3@      L@      @      �?      9@      @     �e@      @      T@      8@                      @     �@@      �?              5@      �?     �^@       @      >@      5@                      @      >@      �?              .@              \@              7@      *@                              @                      @      �?      &@       @      @       @                      ,@      7@       @      �?      @      @      J@      @      I@      @                      $@      .@              �?      @              0@      @      :@      �?                      @       @       @                      @      B@              8@       @              �?      Q@     `e@      &@      0@     �Z@      ,@      |@      8@     �u@      Z@      @              G@      a@       @      "@     �M@      (@      x@      (@     �o@      Q@      @              .@     �D@                      2@      $@     �R@       @      L@      *@      @              ?@     �W@       @      "@     �D@       @     Ps@      $@     �h@     �K@      �?      �?      6@     �A@      @      @      H@       @      P@      (@     �V@      B@              �?      &@      ,@              @      <@       @      >@       @      B@      $@                      &@      5@      @      @      4@              A@      @     �K@      :@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�8hhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?���+@�	           ��@       	                   �2@m[O%+	@�           H�@                           �?��@菛@�            Ps@                           @bpA�&_@R            �_@������������������������       �?����@.            �P@������������������������       �C�Փ�&@$             N@                           @���s`@�            �f@������������������������       ���G�@h            `b@������������������������       �0�<K,@             B@
                           �?���GX�	@*           t�@                          �<@�i%n��@�            �w@������������������������       �*U�F��@�            �s@������������������������       �k����@$            �L@                           @@c��O�	@C           (�@������������������������       �א=�	@�           x�@������������������������       �~��{@(	@K            �]@                           �?i/7c,�@�           �@                          �>@5�?V��@�           ��@                           �?u)�_�@�           �@������������������������       �e��@
           �z@������������������������       ��L�|�?�            `s@������������������������       ��n�x�@             3@                            �?p��i��@�           �@                           @V��9n�@�            0x@������������������������       �2�TF@�            Pu@������������������������       ��Z�@             G@                           @��D�S@�           ��@������������������������       ��!PX��@�            @r@������������������������       ���;���@+           ؊@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        0@     `r@     0�@      ?@     �D@     P}@     �V@     �@     @k@     0�@     pu@      =@      .@     @e@     @l@      6@      :@     �n@      J@      n@     �a@     @p@      i@      5@       @      9@     �F@      @      �?      J@       @      S@      0@     �I@      B@               @      @      2@      @              8@      �?     �B@      @      (@      0@               @       @      "@                      (@      �?      6@      @      @      @                      @      "@      @              (@              .@              @      $@                      3@      ;@              �?      <@      �?     �C@      "@     �C@      4@                      0@      1@                      4@              A@      @      B@      3@                      @      $@              �?       @      �?      @      @      @      �?              *@      b@     �f@      3@      9@      h@      I@     �d@     @_@      j@     �d@      5@      �?      K@      J@       @      @     �J@      @     �N@      ;@     @R@      D@      @      �?      H@      H@       @      @      D@      @     �K@      8@     �P@      9@      @              @      @              @      *@              @      @      @      .@              (@     �V@      `@      1@      2@     `a@     �G@     �Y@     �X@      a@     @_@      2@       @     �S@     �\@      0@      1@      ]@      E@      W@     �R@     �`@     @\@      *@      @      *@      .@      �?      �?      7@      @      &@      8@      @      (@      @      �?      _@     @t@      "@      .@      l@     �C@     ��@     @S@     �@     �a@       @             �C@     @V@              @      H@      @     0u@      .@     �g@      ;@       @             �C@     @V@              @      E@      @      u@      *@     `g@      6@       @              ;@      M@              @     �@@      @     �g@      @      V@      0@                      (@      ?@                      "@              b@      @     �X@      @       @                                              @              @       @      @      @              �?     @U@     `m@      "@      (@      f@      A@     �{@      O@     @v@     �\@      @              ?@     �M@      �?       @      A@      @      a@      4@      S@      7@      �?              <@      K@              �?      A@      �?     �^@      (@     @Q@      2@      �?              @      @      �?      �?              @      *@       @      @      @              �?      K@      f@       @      $@     �a@      >@     `s@      E@     �q@      W@      @              7@      L@      �?      @     �F@      *@      G@      8@      J@      ;@              �?      ?@      ^@      @      @     �X@      1@     �p@      2@     �l@     @P@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJѠ�%hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @=���1@�	           ��@       	                    �?�`A��@p           ��@                           �?�[w�O	@�           Ę@                            �?�P��k@"            |@������������������������       �oHb$C@@�            �m@������������������������       �n@�3��@�            �j@                           �?����	@�           ��@������������������������       �*�I|��@           �z@������������������������       �ZSQ���	@�           �@
                            �?�����*@w           P�@                          �=@�4 �@n            �e@������������������������       ��H�h�@g            �c@������������������������       ��f���/@             .@                           �?<��ZZ�@	           �y@������������������������       �k4J���@h             d@������������������������       ���:�=@�            �o@                           �?yY�-!�@?           8�@                          �5@}_�^�� @i           (�@                           @���?��?�            �y@������������������������       �������?�            �r@������������������������       �"X�����?C            �Z@                           @y�NhϘ@o            �e@������������������������       �>��Q�@9            �V@������������������������       ��ߚ`T@6            �T@                          �7@J���3�@�           $�@                           @�� �@!           ȋ@������������������������       ��k��/�@�            @l@������������������������       ��E'��@�           ��@                            �?o!���@�             q@������������������������       ���`t�@/            @T@������������������������       �fuL�Gj@�            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �r@      �@      =@      K@     Pz@     �Q@     D�@      l@     ȉ@     pu@     �F@      .@     �k@     �s@      6@     �G@     Pr@      I@     @w@     �f@     �w@     �l@     �D@      .@     `e@      o@      4@     �@@     �j@     �A@     �j@     �a@      q@     �f@     �C@      �?      G@     @U@      �?      @      G@      @     @S@      <@     �Y@     �F@      @      �?      <@     �D@      �?      @      2@             �B@      ,@     �O@      7@      @              2@      F@               @      <@      @      D@      ,@     �C@      6@              ,@     @_@     `d@      3@      :@     �d@      >@      a@     @\@     �e@     @a@      @@      @      :@     �Q@      @      *@      O@      @     �R@     �A@     �P@     �L@      "@      &@     �X@      W@      *@      *@      Z@      7@     �O@     �S@     �Z@     @T@      7@              J@     �Q@       @      ,@     @T@      .@     �c@     �C@     �Z@     �F@       @              &@      3@              @      2@      "@     �I@      $@      ;@      2@       @              "@      3@              @      ,@      @     �H@      @      ;@      2@                       @                              @       @       @      @                       @             �D@      J@       @      @     �O@      @     �Z@      =@      T@      ;@                      0@      ,@      �?      @      9@      @     �F@      &@      :@      .@                      9@      C@      �?      @      C@       @      O@      2@      K@      (@                     �S@      l@      @      @      `@      4@     �@      F@     �{@     �\@      @              "@     �Q@      �?      @      ;@      @     �q@      $@      b@      >@                      @     �F@              @      .@             �l@      @      Y@      $@                       @      =@                      &@             �e@      @      T@      @                      �?      0@              @      @              L@              4@      @                      @      :@      �?              (@      @     �J@      @      F@      4@                      @      *@                      @       @     �@@              6@      (@                      �?      *@      �?              "@       @      4@      @      6@       @                     �Q@     @c@      @      @     @Y@      0@     0x@      A@     �r@     @U@      @             �I@     �_@      @      �?     �Q@      ,@     �t@      .@      l@      I@      @              1@     �F@                      .@       @     �U@      @     �@@      *@       @              A@     @T@      @      �?     �K@      @     �n@       @     �g@     �B@      �?              3@      <@      @      @      ?@       @     �K@      3@      S@     �A@      �?              �?      &@                      @              8@      @      :@      (@                      2@      1@      @      @      ;@       @      ?@      0@      I@      7@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJғ�=hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @61��k@�	           ��@       	                    �?��X�O�@|           r�@                           �?����z	@�           @�@                           �?���G�X@4           �}@������������������������       ���h�Ӧ@            @j@������������������������       ������@�            pp@                           �?�aȯ��	@�           ܑ@������������������������       ��rF�G@           �z@������������������������       ����
@�           x�@
                           �?���HL@�           H�@                          �<@�r	��@            �i@������������������������       ��&U>W@v            `g@������������������������       �^�1T\@	             3@                          �4@�iқ#@	           �y@������������������������       �fyp;@|            �i@������������������������       �Ć>1�@�            �i@                           �?|�k�a@*           @�@                          �4@���F@_           ��@                           @09�Xi|�?�            ps@������������������������       ��L����?�            �l@������������������������       �s�H @6            �T@                           �?kb�0	@�             l@������������������������       ��P鷌@P            �_@������������������������       ��Z�@B            �X@                            �?ps@�           ��@                          �:@����?@�           @�@������������������������       �����V�@\           ��@������������������������       �U�O�q�@4            �T@                           @�C���8@;            @������������������������       � y��f@            {@������������������������       �+3Z�@(             P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �s@     ��@      =@      N@     �|@     �R@     ��@     `l@     ��@     �w@      ;@      3@     �k@      t@      3@     �G@     �s@     �J@     pv@      g@     �x@     q@      6@      3@     @f@      m@      .@     �A@     �m@     �C@      l@     �a@     �o@     �k@      3@       @     �C@     �S@      �?      @      P@      �?     �X@      8@     �Z@     �J@      �?       @      ,@      5@                     �@@             �O@      "@     �I@      1@                      9@     �L@      �?      @      ?@      �?      B@      .@      L@      B@      �?      1@     `a@     @c@      ,@      ?@     �e@      C@     @_@      ]@     �b@      e@      2@       @      ;@     �P@       @      "@     �P@      @     �P@      E@     �N@     �Q@      @      .@      \@     �U@      (@      6@     @[@      ?@     �M@     �R@     �U@     �X@      *@             �E@      V@      @      (@      T@      ,@     �`@     �F@     �a@      J@      @              1@      2@               @      *@       @     �R@      @     �N@      (@      �?              .@      .@               @      *@       @     �R@      �?      L@      "@                       @      @                                              @      @      @      �?              :@     �Q@      @      $@     �P@      (@     �N@     �C@      T@      D@       @              @     �D@      @      @      A@             �E@      $@     �C@      7@                      3@      =@              @     �@@      (@      2@      =@     �D@      1@       @      @     �V@     �j@      $@      *@     �a@      5@     ��@      E@      {@     �Z@      @              1@     �N@      �?       @      A@      @     `p@      &@      _@      2@                      (@      8@               @      (@             �f@      @     �P@      @                      $@      4@                      @             @a@      �?      H@      @                       @      @               @      @              F@      @      3@      �?                      @     �B@      �?              6@      @      T@      @     �L@      &@                      @      7@                      0@      @     �J@       @      5@      @                              ,@      �?              @      @      ;@      @      B@       @              @     �R@     @c@      "@      &@      [@      .@     u@      ?@     @s@     @V@      @              H@     �T@       @      @      G@      *@     �g@      :@     �f@     �K@      �?              >@     �Q@       @      @     �A@      *@     �f@      8@      d@     �D@      �?              2@      (@                      &@              @       @      4@      ,@              @      :@     �Q@      @      @      O@       @     �b@      @      `@      A@      @      @      0@      P@      @      @     �H@       @     �`@      @     �]@      @@                      $@      @      @              *@              ,@      �?      $@       @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ� 0hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @����1@�	           ��@       	                    @�-�r�@t           P�@                          �2@Pz���t@�           ,�@                           @�%9�@%           `{@������������������������       �@�� Ƥ@�            �v@������������������������       ��.�Q@.            �Q@                           �?uA� ��@�           T�@������������������������       ��NF��@2           0@������������������������       ����NhZ	@�           ��@
                          �:@��"�� 	@�            �k@                           �?!"3�)@g             e@������������������������       ��PF��
@             @@������������������������       ����G@R             a@                           �?!#+iH	@             J@������������������������       �.��Zz�?             @������������������������       ���w��l@            �F@                          �4@,ְ�@           ��@                           @-ZYUS�@A           ��@                           �?���h@�             l@������������������������       �xؙ�c@B            �Y@������������������������       ��uD/@L            @^@                           �?�ߜR�,@�           ��@������������������������       �T����>�?�             o@������������������������       ��$rkMk@           �{@                           �?z�}�K@�           `�@                           @z�8�@�            �k@������������������������       ���I�׶@#             I@������������������������       �.�Z��@h            `e@                           �?��
{C�@S           x�@������������������������       ��e'3V@�            `o@������������������������       ���xX@�            @s@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     pr@     ��@      .@      J@     �}@     �U@     ��@     `m@     @�@     �t@     �A@      0@      k@     �u@      &@     �D@     �u@     @Q@     �v@     @g@     �v@     �k@     �@@      $@     �g@     `s@      &@     �D@     0s@      L@     �u@     @b@     �u@      j@      4@              1@     �Q@               @      Q@      �?      ^@     �C@     �Q@     �D@      @              (@     �H@              @      P@      �?     @Y@      ?@     �P@     �A@                      @      6@              �?      @              3@       @      @      @      @      $@     �e@     �m@      &@     �@@     �m@     �K@     �l@     �Z@     @q@      e@      1@             �P@     �O@      �?      @     �S@      @     �X@      8@     �[@     �E@      @      $@     �Z@      f@      $@      ;@      d@      I@     ``@     �T@     �d@     @_@      *@      @      <@      B@                     �B@      *@      0@      D@      2@      ,@      *@      �?      8@     �@@                      @@      (@      (@      9@      *@      @      &@              "@       @                      ,@                      �?      @      �?      �?      �?      .@      ?@                      2@      (@      (@      8@      "@      @      $@      @      @      @                      @      �?      @      .@      @       @       @                      �?                                              @      �?       @              @      @       @                      @      �?      @      (@      @      @       @             �S@     �l@      @      &@     �`@      1@     p�@     �H@     �y@     �Z@       @              @@      [@       @      @     �H@      @     �{@      3@     �i@      H@      �?              .@     �D@                      @      @      X@       @     �F@      0@                      $@      2@                      @             �E@       @      2@      "@                      @      7@                       @      @     �J@              ;@      @                      1@     �P@       @      @      F@      �?     �u@      1@      d@      @@      �?               @      3@                      (@             `c@      @      F@      $@      �?              .@      H@       @      @      @@      �?     �g@      &@     @]@      6@                      G@      ^@       @      @     �U@      (@     �j@      >@     �i@     �M@      �?              @      E@                      ,@      $@     �R@      @     �N@       @                      �?      ,@                      @       @      (@      �?      @      @                      @      <@                      $@       @     �O@      @      K@      @                      D@     �S@       @      @      R@       @     @a@      9@      b@     �I@      �?              3@      D@       @      @      B@       @      L@      @     �Q@      3@                      5@      C@              �?      B@             �T@      6@     �R@      @@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJa�>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @*7�U�q@�	           ��@       	                   �1@2����(@�           ҥ@                          �0@��H�g�@#           0~@                           �?�b,:v@a            �c@������������������������       ���1�@            �C@������������������������       �~خ܉�?K            �]@                           @��YW�@�            `t@������������������������       �%���Dq@f            �e@������������������������       ��Kv�A�?\            @c@
                           �?���,j�@�           �@                           �?p�ݖI@�           x�@������������������������       �&i#P�z@�            �p@������������������������       ��n�10�@           P|@                            �?�n�6��@           ܘ@������������������������       ��;�Ƹ@�           X�@������������������������       ��sr�@           z@                           �?��#)�@�           ��@                           �?0�°~@�            Pv@                           �?u�<S�)@�            �i@������������������������       �����@A            �X@������������������������       �{�0���@@            �Z@                           @(q���?Y             c@������������������������       ��]Jgnc@            �G@������������������������       �ڝ��8��?>            �Z@                           @��â	@�           ؇@                           @��ch^	@p            �@������������������������       �R����@�            �x@������������������������       �K� ��[	@{             g@                          �3@�!d7v@y            `g@������������������������       �����KK @*            @P@������������������������       �/���"@O            �^@�t�b�~     h�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     (�@      C@     �Q@     �y@     �T@     �@     �k@     �@     �v@      @@      &@      l@     �w@      2@     �G@     `q@     @P@      �@     �c@     0�@     �m@      5@      �?      2@     �P@              @      @@      @      k@      *@     �X@      =@                      @      >@                      ,@              R@      �?      6@      *@                      @      @                      "@              "@              @      @                      �?      7@                      @             �O@      �?      2@      @              �?      *@      B@              @      2@      @      b@      (@     @S@      0@              �?      @      9@                      *@      @     �N@       @      C@      0@                      @      &@              @      @              U@      @     �C@                      $@     �i@     �s@      2@      E@     �n@      O@     8�@     @b@     0~@     @j@      5@              N@     �X@      @      @      N@      &@      n@      >@     �c@      J@      �?              >@      A@       @      @     �@@       @      I@      3@      K@      B@      �?              >@     @P@      �?      �?      ;@      "@     �g@      &@     �Y@      0@              $@     `b@     �j@      .@      B@     @g@     �I@     ps@      ]@     `t@     �c@      4@       @      \@     �d@      $@      ?@     �]@     �C@     �k@     @X@     @o@      Z@      1@       @     �A@      I@      @      @     �P@      (@     @V@      3@      S@      K@      @      "@     �R@      e@      4@      7@     @`@      2@     `p@      O@     `k@     �^@      &@              6@      I@       @      @     �A@             `a@      2@      Q@      4@                      ,@     �D@       @      @      ;@             �J@      ,@      @@      2@                      @      ,@       @       @      2@              <@      @      1@      @                      "@      ;@              �?      "@              9@       @      .@      (@                       @      "@                       @             �U@      @      B@       @                      @      �?                      @              4@      @      *@      �?                      @       @                      @             �P@              7@      �?              "@      J@     �]@      2@      4@     �W@      2@     �^@      F@     �b@     �Y@      &@      "@     �F@     @Y@      $@      0@     @T@      1@      P@      E@     �W@     @V@       @      @      >@     �O@       @      &@     @P@      *@      C@      .@     �Q@     @Q@      @      @      .@      C@       @      @      0@      @      :@      ;@      7@      4@      @              @      2@       @      @      ,@      �?     �M@       @     �L@      ,@      @               @      $@                      @              5@      �?      9@                              @       @       @      @       @      �?      C@      �?      @@      ,@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�k�\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @~�uNi�@�	           ��@       	                    �?XzU,ގ@�           ��@                          �<@�eY9'@�           ��@                          �1@�w%d@�           ؃@������������������������       �Z!�� @A            �Y@������������������������       �vIg��@S           ��@                          �?@�?�7�1@)             Q@������������������������       �)���@             H@������������������������       ��6,؊� @
             4@
                          �1@�i��e6	@�           X�@                          �0@��n�$�@q            @f@������������������������       ��ڙ��@             �L@������������������������       �#�M��@Q            @^@                           �?�����o	@a           ��@������������������������       �U��[��@�            �w@������������������������       �3�Iw��	@o           (�@                           �?�G�=E@           Й@                            �?i��&� @]           (�@                           �?��R�W�?M             _@������������������������       �c3`o���?(            @P@������������������������       �-�x.��?%            �M@                          �5@���&@           �z@������������������������       ��勑u� @�            s@������������������������       ���]�� @P             ^@                           @�r�op.@�           <�@                          �<@/��S�@�           Є@������������������������       ��Λ��Q@�           �@������������������������       �E�t��r@             =@                          �5@��&V@           P{@������������������������       ��2P��@�             p@������������������������       �l�BC�@p            `f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        @      r@      �@     �@@      N@     P|@     @R@     �@     @j@     �@     Pt@      ;@      @     @j@     0t@      8@     �G@     �s@      O@     �z@      g@     �y@      m@      8@             �N@      W@      �?      (@     @U@      @     `h@      B@      d@     �H@      @              K@     �T@      �?      "@      S@      @     @h@      ;@     �b@     �@@       @               @      *@                      $@              H@      @      7@      @                      J@     �Q@      �?      "@     �P@      @     @b@      8@     �_@      =@       @              @      "@              @      "@              �?      "@      &@      0@      @               @      @               @       @              �?      "@      @      0@      @              @       @              �?      @                              @                      @     �b@     �l@      7@     �A@     �l@      L@     �l@     �b@      o@     �f@      3@      �?      "@      A@               @      .@             �F@      .@      D@      1@                      @      .@               @      "@              ,@      �?      @      @              �?      @      3@                      @              ?@      ,@     �@@      &@              @     �a@     �h@      7@     �@@     �j@      L@      g@     �`@      j@     �d@      3@              9@     �Q@       @      *@      N@      @     �L@      F@     �K@     �E@      @      @     �\@     �_@      5@      4@     `c@     �H@     �_@     @V@      c@     �^@      (@              T@     �k@      "@      *@     @a@      &@     Ȅ@      :@     �x@     @W@      @              *@     �Q@      @       @      @@      @     �p@      @      `@      1@      �?                      "@      @              @      @     @T@      �?      0@      @                              @                       @             �F@              $@      @                              @      @              @      @      B@      �?      @      �?                      *@     �N@               @      :@       @     �g@      @     @\@      (@      �?              &@     �C@               @      3@       @     �b@      @     @R@      @      �?               @      6@                      @             �D@              D@       @                     �P@     �b@      @      &@     �Z@      @     �x@      4@     �p@      S@       @              7@     @Z@      @      $@      N@      @     �l@      (@      f@     �F@                      3@     �Y@      @      $@      I@      @     `l@      &@     �e@      C@                      @      @                      $@              �?      �?      @      @                      F@      G@      @      �?      G@      @     �d@       @     �U@      ?@       @              2@      =@              �?      $@      @      ^@      �?     �M@      0@      �?              :@      1@      @              B@              G@      @      <@      .@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJc7(hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @n��}T@�	           ��@       	                    �?��)[ 	@s           .�@                            �?r�8@�Y@�           x�@                           �?��&ܚ�@�            �h@������������������������       �ը~�7�@_            `a@������������������������       �ӫA��@&            �L@                          �<@�4Oa@           �|@������������������������       �
���@�            `y@������������������������       � �֌mm@"            �J@
                          �9@hP�w٭	@�            �@                           �?�>�(0	@�           l�@������������������������       �}���	@           ��@������������������������       ��3��@�            Pt@                           @����t�
@�            �v@������������������������       ��f��u�
@�             s@������������������������       � ��@$            �N@                          �1@�+��D�@D           Ț@                           @xX��u�?�            �w@                           �?T�q;��?8            �V@������������������������       �&r�1a�?            �F@������������������������       �fT����?            �F@                          �0@P,�4���?�            Pr@������������������������       �"\.<�c�?<            �Y@������������������������       �pbF�H�?q            �g@                          �8@��pU�@_           ̔@                           @(�p]�@�           ��@������������������������       �fsÇ��@�             n@������������������������       �����p@�           (�@                           �?�ܕˇ�@�            �s@������������������������       ����S�@W            �a@������������������������       �N U�RK@q             f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@      r@     x�@      @@     �L@     @}@      U@     �@      n@     ��@     @u@      <@      4@     �i@     s@      :@     �G@      t@      O@     �w@      i@     �w@     @l@      :@              L@     �U@      @      $@     �U@      @     �c@      ?@     �c@     �M@       @              .@      :@              @      7@      @     �C@      @     @P@      *@      �?              ,@      1@              �?      3@       @      9@      @     �E@      &@      �?              �?      "@              @      @      �?      ,@              6@       @                     �D@     �N@      @      @      P@       @     �]@      9@      W@      G@      �?              C@     �K@      @      @      K@       @     �\@      0@     �V@      >@      �?              @      @               @      $@              @      "@       @      0@              4@     �b@     @k@      7@     �B@     `m@     �L@     �k@     @e@     �k@     �d@      8@      *@     �Z@     �f@      .@      :@     �h@      <@     �g@     �\@     `g@     �Z@      .@      *@     �T@     �]@      .@      5@     @b@      5@      \@     @W@     �`@     �T@      .@              8@     �N@              @      J@      @     @S@      6@      J@      9@              @      F@      C@       @      &@     �B@      =@      A@     �K@     �@@      N@      "@       @      D@      A@      @      &@      ?@      ;@      ?@      ?@      >@     �I@      "@      @      @      @      �?              @       @      @      8@      @      "@                      U@     �k@      @      $@     @b@      6@     P�@     �C@     0z@     �\@       @              @     �C@              �?      4@             �j@       @     �U@      1@                      �?      &@                      �?             �K@              ,@       @                      �?      @                      �?              8@              @       @                              @                                      ?@              $@                              @      <@              �?      3@             �c@       @      R@      "@                      �?      2@                      @              J@              1@       @                       @      $@              �?      *@             �Z@       @     �K@      �?                      T@     �f@      @      "@     �_@      6@     @{@     �B@     �t@     @X@       @              N@      a@      @      @     �U@      0@      w@      .@     �o@     �P@       @              3@      E@       @              3@      $@     �Q@      @     �O@      (@      �?             �D@     �W@       @      @     �P@      @     �r@      (@     �g@     �K@      �?              4@      G@       @      @      D@      @     �P@      6@     @T@      >@                       @      7@               @      ,@              E@      @     �@@      *@                      (@      7@       @       @      :@      @      8@      0@      H@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?BB?�CC@�	           ��@       	                   �8@�����P	@�           ��@                          �1@5���@�           ��@                           �?�M�Q��@{            �g@������������������������       �"�H��`@1            �R@������������������������       �^r��Z@J            �\@                           �?�;BǏ	@H           X�@������������������������       �&��L�d@�             v@������������������������       �{���#+	@i           H�@
                          �:@#���>�	@;           p@                           �?�0v��s@n            �d@������������������������       ��T��-@%             M@������������������������       �l�}�y�	@I            @[@                           �?+|�׮	@�             u@������������������������       �\L�L�D@:            �Y@������������������������       �0c���w	@�            @m@                            �? ;� &�@�           ҡ@                          �4@L��;��@9           �@                           @%*I=��@�           x�@������������������������       ��f�j�N@l            �f@������������������������       �ϯ��:�@P           ؀@                          @@@\3�<�@}           P�@������������������������       �l8��9V@u           ؂@������������������������       �ɮ<
�@             .@                            @�scЊ.@k           ��@                          �7@W����@X           �@������������������������       �tn�>�@           �x@������������������������       ��z��V�@Q            �^@                          �9@�{�Y��@           �z@������������������������       ����FV�@�             v@������������������������       �Vl��q+@6             S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@      �@      9@     �M@     p{@     @T@     ��@     �j@     ��@     @v@     �B@      1@     �d@     @o@      .@     �E@      o@     �E@      l@     �a@     �o@     �i@      >@      $@     �]@     @d@      (@      ;@      f@      3@     �f@     @T@     �i@      ^@      .@              (@      @@      �?      �?      5@      �?     �J@      (@      E@      .@                              ,@      �?              @      �?      9@      @      (@      "@                      (@      2@              �?      ,@              <@      @      >@      @              $@     �Z@     @`@      &@      :@     �c@      2@     @`@     @Q@     `d@     @Z@      .@      @      8@     �P@       @      .@      K@      @      K@      2@     �Q@     �A@      @      @     �T@      P@      "@      &@     �Y@      (@      S@     �I@      W@     �Q@      "@      @     �G@      V@      @      0@     �Q@      8@     �D@     �M@     �G@     @U@      .@              1@     �F@       @      @      1@      @      .@      5@      3@      1@       @              "@      6@                      @              @      @       @      @                       @      7@       @      @      *@      @      $@      0@      &@      (@       @      @      >@     �E@      �?      *@      K@      5@      :@      C@      <@      Q@      @               @      1@              @      2@      �?      3@      @      &@      1@              @      6@      :@      �?      @      B@      4@      @     �@@      1@     �I@      @       @      `@     `r@      $@      0@     �g@      C@     ��@     �R@     Ё@     �b@      @              V@     �f@      @      $@      [@      >@     �{@     �D@     @u@     �T@      @              C@     @V@      @      @     �K@      @     r@      *@     �f@     �E@                      &@      @@      �?       @      4@      @     �J@      @     �D@      (@                      ;@     �L@       @       @     �A@             �m@       @     �a@      ?@                      I@     �W@       @      @     �J@      ;@     �c@      <@     �c@     �C@      @             �H@     @V@       @      @     �J@      6@     �c@      :@     �c@      C@      @              �?      @                              @               @      �?      �?               @      D@     �[@      @      @     �T@       @      v@      A@     �l@     @Q@       @       @      1@      N@      �?      @     �H@      @     `i@      .@      `@      <@       @              0@     �I@      �?      @      >@      @      f@       @     @U@      .@       @       @      �?      "@                      3@      �?      ;@      @     �E@      *@                      7@     �I@      @      @      A@       @     �b@      3@     �Y@     �D@                      3@      G@      @              9@       @     @`@      $@      U@     �A@                      @      @      �?      @      "@              5@      "@      2@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�"�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�G?Ru@�	           ��@       	                    �?#(BD�@a           .�@                           �?�5��"@�           ��@                           �?�%��6P@�            �m@������������������������       ��UO;@��?A            �X@������������������������       ����n
@Z             a@                            �?�"AN��@C            �@������������������������       ��o����@f            �b@������������������������       �˵���	@�            �v@
                           @�L���v@�           ��@                           �?��t��g@�            �u@������������������������       �&����@I            �\@������������������������       ��q��Q�@�             m@                            �?�S[�@�           ,�@������������������������       ������?�            �m@������������������������       �)5�@           ��@                           �?�YA�	@?           Ț@                           �?6�b�M
@&           0�@                            @f�A`�	@�             u@������������������������       ������@s             g@������������������������       �Wbm$�j
@e             c@                           �?�@]u
@N           ��@������������������������       ��ؿW��@M            @_@������������������������       �bʟ���
@           py@                           �?!�f|/�@           `�@                          �=@�e���u@�            `k@������������������������       �-�-�@y            `h@������������������������       ��Jz��@             8@                           @m�I�W@�           ��@������������������������       ���9�@q             g@������������������������       ��K?�@!           �{@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@      r@     @�@      ;@      P@     P}@      V@     h�@     �k@     ��@     �u@     �@@      @      ]@     �s@      @      ?@      m@     �@@     8�@     @W@     �~@     @c@      &@      @     @P@     @Y@      @      2@      `@      ,@     �`@      K@      c@     @Q@      @              1@      B@              @      7@      �?      Q@      0@      L@      0@                              3@                       @             �B@       @      @@      �?                      1@      1@              @      .@      �?      ?@      ,@      8@      .@              @      H@     @P@      @      .@     �Z@      *@     �P@      C@      X@     �J@      @              1@      1@                      ?@      �?      8@      0@      <@      (@      @      @      ?@      H@      @      .@     �R@      (@      E@      6@      Q@     �D@       @             �I@     �j@      �?      *@      Z@      3@     �@     �C@     @u@     @U@      @              $@     �L@      �?      @     �@@      @      \@      9@     @Q@      >@                      @      @               @      $@       @     �F@       @     �@@      $@                      @     �I@      �?       @      7@      @     �P@      7@      B@      4@                     �D@     `c@              "@     �Q@      (@     }@      ,@     �p@     �K@      @              @      7@               @      ,@             @_@       @     �J@      .@                      C@     �`@              @     �L@      (@     @u@      (@     @k@      D@      @      2@     �e@     �m@      5@     �@@     �m@     �K@     `r@     @`@     �r@     @h@      6@      2@      X@      `@      0@      ;@      _@      C@      W@     @T@     �]@     �[@      3@      @      @@     �K@      @      @      J@      .@     �D@      C@     �@@      I@       @      �?      2@      =@                      ?@      $@      :@      <@      *@      ;@       @      @      ,@      :@      @      @      5@      @      .@      $@      4@      7@      @      (@      P@     �R@      &@      8@      R@      7@     �I@     �E@     �U@     �N@      &@              ,@      9@                      2@              3@      @      9@      ,@      @      (@      I@     �H@      &@      8@      K@      7@      @@     �C@     �N@     �G@      @             �S@     �[@      @      @      \@      1@     @i@     �H@     `f@     �T@      @              *@      <@                      5@      @     �T@      @      F@      2@      �?              (@      <@                      2@      @     @S@      �?     �D@      .@                      �?                              @      @      @      @      @      @      �?             @P@     �T@      @      @     �V@      &@      ^@     �E@     �`@     @P@       @              7@      @@              @      7@      @      6@      9@      @@      2@      �?              E@      I@      @      @      Q@      @     �X@      2@     �Y@     �G@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJM2�1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?%,�v@�	           ��@       	                    �?,�%�M�@           ��@                           �??x?7I�@>           @                            @���<7@v            @g@������������������������       �ƞyO�#@Z            �a@������������������������       �!��O� @            �F@                          �<@�=gf$@�            ps@������������������������       ��?6lA�@�            �p@������������������������       �X�M� x@            �E@
                            �?	�L�@�           ��@                           �?�?�1f@z            �j@������������������������       ��gm��?=            �Z@������������������������       �誱�@=            �Z@                            @���o�@\           �@������������������������       ��|��W@           �y@������������������������       �0��ooS�?U            �`@                          �5@1ʢ<d@�           ¤@                          �1@s��T�@i           ��@                           @LvA�t@�            0v@������������������������       ��U�=�@%             I@������������������������       �����>I@�            s@                           �?wsE�o@�           �@������������������������       �v
[�@1             T@������������������������       ���MB\@T           ��@                           @� ��U	@,           �@                          �;@6|��b�	@           ��@������������������������       �$����e	@y           0�@������������������������       ��O�
@�            @m@                           @���9�@           �|@������������������������       �<3ע�1@�            �s@������������������������       ������j@b            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �t@     ȁ@     �@@     �J@     �z@      V@     Ȏ@      k@     ��@     �x@      @@      @     �V@      g@      @      @      V@      $@     �{@      E@     0r@     @W@      @      @     �O@     @T@      �?      @      H@       @      W@      >@     @]@      J@      @      @      *@      5@                      1@              G@      @      L@      5@      �?      @      (@      .@                      0@              >@      @      C@      3@      �?              �?      @                      �?              0@      �?      2@       @                      I@      N@      �?      @      ?@       @      G@      7@     �N@      ?@       @             �G@      J@      �?       @      :@       @      F@      4@     �K@      1@       @              @       @               @      @               @      @      @      ,@                      ;@      Z@       @      �?      D@       @     �u@      (@     �e@     �D@       @               @      >@       @              ,@      @     @Z@             �C@      .@       @                       @                      @       @      P@              .@      (@                       @      6@       @              "@       @     �D@              8@      @       @              9@     �R@              �?      :@      @     `n@      (@     �`@      :@                      2@     �P@                      3@      @      e@      $@     �Y@      9@                      @      @              �?      @             �R@       @     �@@      �?              "@     �n@      x@      >@      H@      u@     �S@     �@     �e@     �}@      s@      ;@       @     �W@     �j@       @      0@     `a@     �@@     �w@     �N@     �q@     �a@      .@              3@     �I@              @      =@       @     �]@      *@     @V@      :@                      @       @                      @              9@      @      @      @                      ,@     �H@              @      :@       @     �W@       @     @U@      4@               @     �R@      d@       @      "@     �[@      ?@     p@      H@     �h@     �\@      .@              @      :@              �?      ,@      @      @      @      *@      "@               @     �Q@     �`@       @       @      X@      ;@     `o@     �F@     �f@     @Z@      .@      @     �b@     �e@      6@      @@     �h@     �F@      e@     @\@     �g@     �d@      (@      @     �W@     �Z@      2@      ;@     @`@     �C@     �Q@     �V@      Y@     �^@      (@      �?     �P@     �R@      "@      3@      Y@      3@     �N@     �P@     �T@     @R@      "@      @      ;@     �@@      "@       @      >@      4@      $@      7@      1@     �H@      @      �?      L@     @P@      @      @     �P@      @     �X@      7@     �V@      F@              �?      @@     �G@              �?      H@      �?     @V@      "@      N@      8@                      8@      2@      @      @      3@      @      "@      ,@      ?@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@/�v,9@�	           ��@       	                    @�;>�J@�           |�@                           @�;�@�           ��@                           �?ܽ�>!@]           �@������������������������       ���2��@u            @g@������������������������       ��Mj�@�            �v@                           @np:J�=@[             b@������������������������       ����1s�@=            �X@������������������������       �ŕ�>�@            �F@
                           @M����� @�           `�@                           �?H��� @�           h�@������������������������       ����W(�?�            Pr@������������������������       ���`��@
           �z@                            �?.A�%� @             ?@������������������������       ��8��jZ�?             7@������������������������       �      �?              @                           �?���;�h@&           T�@                           �?��s�l�@�           X�@                           �?.�=��4@�            pt@������������������������       �yVǎd@O            �a@������������������������       �r���#x@n             g@                            �?y�y�@�            @x@������������������������       ��R�`I@6            �S@������������������������       ����6@�            Ps@                           @���~	@u           |�@                           @I�8A�@�           �@������������������������       �j 
b�Z	@d           ��@������������������������       ���j^�[@z           ��@                           �?�C�Ҧ�	@�            �l@������������������������       ����4�	@>            �W@������������������������       �}���@Y            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �r@     p�@     �C@     �H@      ~@     �L@     (�@      i@     �@     �t@      F@      @      R@      g@      @      @      a@       @     �@     �J@     �v@     �W@      @      @     �L@     �V@      @      @      X@      @     �c@     �E@     @d@     �P@      @       @     �C@     �N@      @      @     �S@      @     �^@     �@@     `b@      K@                      @      <@      @              G@      �?     �C@      ,@      A@      ,@               @      @@     �@@      �?      @      @@      @     �T@      3@     @\@      D@               @      2@      =@                      2@       @     �A@      $@      .@      (@      @      �?      2@      6@                      @              9@      @      @      (@       @      �?              @                      &@       @      $@      @       @              �?              .@     �W@      @      @      D@       @     v@      $@     �h@      =@                      ,@     �V@      @       @      C@       @     u@      $@     �h@      7@                      @      @@              �?      "@              d@      @     �R@      @                       @     �M@      @      �?      =@       @      f@      @     �^@      0@                      �?      @              �?       @              0@               @      @                              @              �?      �?              (@                      @                      �?                              �?              @               @                      0@     `l@     `w@      @@     �E@     �u@     �H@     p~@     `b@     �}@      n@     �D@      �?      N@     �W@       @       @     �R@      @     `j@      <@     �e@      G@      $@      �?      H@      H@      �?      @      C@             �I@      .@      T@      ?@      "@      �?      5@      2@                      1@             �B@      @     �A@      @      @              ;@      >@      �?      @      5@              ,@      (@     �F@      8@      @              (@     �G@      �?      @     �B@      @      d@      *@     �W@      .@      �?                      "@      �?      �?      ,@       @      =@      �?      ,@      @      �?              (@      C@               @      7@       @     ``@      (@     @T@       @              .@     �d@     pq@      >@     �A@     �p@     �F@     @q@     �]@     �r@     @h@      ?@      "@      a@     �m@      ;@     �@@      n@      E@     �n@      W@     @q@     �e@      0@      @     �X@     �d@      9@      7@     �e@      ?@     �X@      R@     �_@     �^@      ,@      @     �B@     @R@       @      $@     �P@      &@     `b@      4@     �b@     �I@       @      @      ?@      D@      @       @      >@      @      >@      ;@      5@      5@      .@      @      @      2@      �?              .@      �?      $@      ,@      @      &@       @              8@      6@       @       @      .@       @      4@      *@      2@      $@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��ShG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                            �6@P�[�h@�	           ��@       	                    @���),5@'           (�@                           �?�Gg���@�           �@                           �?���8��@G           P@������������������������       �D���E<@�            �m@������������������������       ��,��Y�@�            pp@                          �3@.���o�@�           @�@������������������������       �o:�*�t@d           �@������������������������       ���6�D	@5           �~@
                           @�}]��(@G           x�@                           �?�����4 @�            �@������������������������       �����r��?�             j@������������������������       ��6���~@�            0y@                            �?��=��@�            �r@������������������������       �[V��@'             N@������������������������       �VBl��h@�            �m@                          �<@�[��@�           Ԗ@                           �?[y�5/@�           ��@                           @ۊ�[	@H           0�@������������������������       ����>@�            @n@������������������������       �p`���	@�            @q@                           @pOv1;w@           ؂@������������������������       �����@           �{@������������������������       �����@d            `d@                          �A@K��T	@�            @u@                            �?+�U�w�@�            �t@������������������������       ���0۸@q            �g@������������������������       �
H+z�`	@\            `a@������������������������       ��+��>3�?             (@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        4@     Ps@     `�@      ?@     �H@     �}@     @T@     P�@      n@     ��@      w@      8@      $@      e@      w@      (@      9@      p@      C@     `�@      `@     �@     �f@      &@      $@     �a@      m@      $@      0@      g@      B@     `u@     @]@     `s@     @`@      $@              E@      T@              �?     �F@      @     �c@      8@      ]@      >@      �?              3@     �A@              �?      5@      @     �U@      1@      D@      *@      �?              7@     �F@                      8@             �Q@      @      S@      1@              $@     @Y@      c@      $@      .@     `a@      ?@      g@     @W@     @h@      Y@      "@      @     �D@     �S@              @     �Q@      &@      `@     �I@     �V@     �N@      @      @      N@     �R@      $@      &@      Q@      4@      L@      E@      Z@     �C@      @              :@     �`@       @      "@      R@       @     `y@      &@     @h@     �J@      �?              $@     @V@              @      A@             `s@      @      `@      ?@                      @      <@                      @             @`@             �B@      @                      @     �N@              @      ;@             �f@      @      W@      ;@                      0@      G@       @      @      C@       @      X@      @     @P@      6@      �?              @      @                       @              :@              &@      @                      $@     �E@       @      @      >@       @     �Q@      @      K@      0@      �?      $@     �a@     �g@      3@      8@     �k@     �E@     �k@      \@     �q@      g@      *@      @      Z@     @c@      (@      2@     �e@      :@      h@     @S@     `m@      \@      &@      @      N@     @R@      "@      &@     �U@      1@      J@      H@     @V@     �M@      $@      �?     �B@      >@      �?      @     �D@      @      6@      1@     �L@      3@      @       @      7@     �E@       @      @      G@      &@      >@      ?@      @@      D@      @      �?      F@     @T@      @      @      V@      "@     �a@      =@     @b@     �J@      �?      �?      A@     �L@               @      N@      @     �\@      2@     �Y@     �F@      �?              $@      8@      @      @      <@      @      :@      &@      F@       @              @      B@      A@      @      @      H@      1@      =@     �A@     �G@     @R@       @      �?      B@      ?@      @      @      H@      1@      =@     �A@      G@     �Q@       @              5@      3@               @      7@      *@      (@      3@      =@     �H@       @      �?      .@      (@      @      @      9@      @      1@      0@      1@      5@              @              @                                                      �?      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJa�fhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                              @�T�6�!@�	           ��@       	                     �?���7�@�           ��@                           @G���@?           ��@                           �?�P�}
�@�           ��@������������������������       ����Q[@�            �w@������������������������       ��\ٰx	@�           ��@                            �?U�,���@`           H�@������������������������       �݂�gF@�             y@������������������������       ��#q}�@f           ��@
                           �?�����@�           ��@                           @"�EG�@�            �s@������������������������       ��ꀁ��@B            @Y@������������������������       �F�3|�a@�            `j@                          �:@�T��>�@�            �u@������������������������       �.� 8�#@�            �r@������������������������       ��lB ;@             G@                           @W�Z�@�           ȑ@                           �?P��D{�@           P�@                           �?u��H	@�            u@������������������������       �`����f@F            @\@������������������������       �z#�N�	@�             l@                          �4@�5?�Ss@;           �@������������������������       �z�Lt�s@�            @k@������������������������       ��w/ƥ@�            �q@                           @y���L�@�            �r@                          �9@��+ee @Q            �`@������������������������       �aY[Y��?G            @]@������������������������       ��1H����?
             0@                           �?�D����@^            `d@������������������������       �뛩�\�@*            @R@������������������������       �39&��@4            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        8@     0s@     ��@      7@      I@     �|@     @T@     ؏@     @i@     ��@     �t@      =@       @     `i@     0y@      *@     �@@     0s@      J@     x�@     �a@     0�@     �l@      4@      @      c@     �s@      &@      =@     �j@      D@     �@      \@     ~@      h@      0@      @     �Z@     �d@      "@      :@     �a@      @@     @k@     �U@     @l@     @]@      ,@      �?      =@      H@              @      A@      �?     �Z@      0@     �Z@      @@      @      @     @S@      ]@      "@      5@     @[@      ?@     �[@     �Q@      ^@     @U@      &@              G@      c@       @      @     �Q@       @     �t@      9@     �o@      S@       @              4@     �H@              �?      8@             �e@      &@     �V@      ?@                      :@      Z@       @       @     �G@       @      c@      ,@     �d@     �F@       @      �?     �I@     �U@       @      @     @W@      (@     �i@      =@     �`@     �B@      @      �?      7@     �C@      �?      �?      F@      @     �X@      *@      M@      ;@       @      �?      &@      "@                      2@      @      *@      $@      2@      1@                      (@      >@      �?      �?      :@             �U@      @      D@      $@       @              <@     �G@      �?      @     �H@       @     �Z@      0@     �R@      $@       @              6@     �F@              @      <@      @      Y@      .@     �P@      $@       @              @       @      �?              5@      �?      @      �?       @                      0@      Z@      d@      $@      1@     �c@      =@     �p@     �N@     @j@     �X@      "@      0@     @V@     �`@      "@      (@     �`@      ;@      b@     �L@      a@     �S@      "@       @      =@     �J@      @      @     �J@      2@      M@      ,@     �J@     �A@       @              &@      .@              @      3@      �?      =@      @      4@      $@               @      2@      C@      @      @      A@      1@      =@      "@     �@@      9@       @       @      N@     �S@       @      @     �S@      "@     �U@     �E@     �T@      F@      @      @      ,@      9@              @      >@       @     �K@      0@      H@      ,@      @      �?      G@      K@       @      �?     �H@      @      ?@      ;@     �A@      >@      @              .@      <@      �?      @      8@       @      _@      @     �R@      3@                      @       @              @      @      �?      S@      @      9@      @                      @       @              �?      @      �?     �Q@      �?      5@      @                                              @                      @      @      @                              $@      4@      �?      �?      3@      �?      H@             �H@      ,@                              (@                       @      �?      5@              8@      @                      $@       @      �?      �?      &@              ;@              9@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJT�V3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?(�O�g@�	           ��@       	                    �?p�/6|@�           p�@                           �?*h5<�U@(           �}@                          �1@O��@r            @e@������������������������       ��
ڬu��?             :@������������������������       ��t;c@b             b@                          �7@/dQY@�             s@������������������������       �X91�@v            @h@������������������������       ������d@@            �[@
                          �2@��5@�           �@                            �?��ż-�?�            �q@������������������������       �86u�*�?3            �T@������������������������       �<�E�&& @�            `i@                           @��A2(@           @z@������������������������       �LG�+��@~            �i@������������������������       ��L.Q�� @�            �j@                           @<��M@�           Z�@                           @�M��@�           ܢ@                           �?H�F�Yp	@�           @�@������������������������       �'9 ���	@U             b@������������������������       �'�fw�7	@+           ��@                           �?~���o@}           ��@������������������������       ��3��Q@4            @U@������������������������       ��>��0�@I           H�@                            �?܊��G	@�            �s@                            �?��~	@p            �f@������������������������       �գ�ʆ;@9            �W@������������������������       ��tm��/@7            @U@                           �?JuE��@X            `a@������������������������       ����g�@!            �I@������������������������       ���u?�@7             V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     ��@     �@@     �R@     0~@     @S@     ��@      i@     ��@     Pu@      8@              U@      d@      @      ,@     @Y@      @     `z@     �B@     �p@     �S@      @             �M@     �Q@       @      ,@      L@      @     �V@      8@     @Y@      I@      @              0@      7@                      0@              F@      @      J@      ,@                       @                              @              (@               @                              ,@      7@                      (@              @@      @      F@      ,@                     �E@      H@       @      ,@      D@      @     �G@      3@     �H@      B@      @              ?@      ;@       @      @      6@      �?     �E@       @      B@      4@      �?              (@      5@              &@      2@       @      @      &@      *@      0@       @              9@     �V@      �?             �F@      @     �t@      *@      e@      =@                       @      ;@                      0@             �c@              N@      1@                              "@                      @             �M@              "@       @                       @      2@                      (@             �X@             �I@      .@                      1@     �O@      �?              =@      @     �e@      *@     @[@      (@                      *@      2@                      2@      @     @T@      @      M@      @                      @     �F@      �?              &@              W@      @     �I@      @              9@     �l@     Pw@      >@     �N@     �w@     �Q@     P�@     �d@     ��@     `p@      5@      0@     �h@     �t@      <@      M@     �u@     �N@     H�@      _@      ~@      m@      *@      .@     @a@      h@      9@      F@      o@     �K@      j@     �Y@     �j@     @e@      *@      @      0@      (@              (@     �@@      @      "@      ,@      2@      1@      @      $@     �^@     �f@      9@      @@     �j@     �H@     �h@      V@     `h@      c@      $@      �?      M@     �a@      @      ,@     @Y@      @     �s@      6@     �p@     �O@              �?      @      4@              �?       @      @      ,@      @      7@      @                      K@     �^@      @      *@     @W@             �r@      3@     �n@      M@              "@     �@@      C@       @      @     �@@      $@     @P@      D@     �H@      =@       @      @      5@      0@       @       @      $@       @      C@      =@      =@      1@       @              *@      &@       @      �?      @       @      0@      ,@      0@      ,@      �?      @       @      @              �?      @      @      6@      .@      *@      @      �?      @      (@      6@              �?      7@       @      ;@      &@      4@      (@      @      @              &@              �?       @       @      $@      @      @      @       @              (@      &@                      .@              1@      @      1@      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�G�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���Bc@�	           ��@       	                   �1@�8�U�@@r           ��@                           @�H6m�W@�           ��@                           @_����� @�            r@������������������������       �d
�@Q             \@������������������������       �n��E�T�?j             f@                           �?mSo�'@�            �s@������������������������       ��a�@5            �S@������������������������       ���m�-@�            �m@
                           �?pD�8_@�           ��@                           �?�ø/j�@           0z@������������������������       �(�oG
@[            `a@������������������������       �E�?l@�            �q@                          �3@�E�=@�           �@������������������������       �Q#Tu5@>            �@������������������������       �$G)9@�             o@                            @�~~O�@6           ��@                           @����@�           ��@                           @&hŎ�e	@�           @�@������������������������       �S�V�
"	@�           P�@������������������������       �����=@9            �W@                          �5@i�}ߗ-@�           ��@������������������������       �f��l�Z@`            �b@������������������������       �����v@M           0�@                           �?U�I��@�           0�@                           @�顩��@�            �n@������������������������       �QIU��Q	@�            �g@������������������������       ��7a[+�@$            �K@                          �:@��V�@�            w@������������������������       ��!�Mo.@�            �m@������������������������       �'�@N            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     H�@      B@      M@     �|@     @R@     <�@      m@     �@      w@      B@       @     �T@      m@      (@      $@     `e@      3@     Ѓ@     �T@     �w@     @b@      &@      �?      1@     �R@      �?      @      E@             pq@      9@      `@      @@       @               @      :@              @      ,@             @d@      ,@     �G@      *@       @              @      $@                      $@              H@      (@      4@      @                      @      0@              @      @             �\@       @      ;@      @       @      �?      "@     �H@      �?      �?      <@             @]@      &@     �T@      3@              �?      @      &@      �?              .@              0@       @      0@      (@                      @      C@              �?      *@             @Y@      "@     �P@      @              @     �P@     �c@      &@      @      `@      3@     0v@      M@     �o@     �\@      "@      @      @@     �F@      @       @      O@      *@      R@     �C@     @T@      J@      "@      @      $@      7@      �?      �?      =@      @      <@      2@      $@      &@      �?      @      6@      6@      @      �?     �@@      $@      F@      5@     �Q@     �D@       @              A@      \@      @      @     �P@      @     �q@      3@     �e@      O@                      5@     �R@       @      �?     �F@       @     �g@      &@     �`@      B@                      *@     �B@      @      @      6@      @     �W@       @      C@      :@              "@      k@     r@      8@      H@     r@      K@     Py@     �b@     Px@      l@      9@      @      c@     �h@      *@      B@     @k@     �E@      r@     @X@     `r@     �a@      3@      @     �[@     �Y@      "@      ;@      `@      7@      [@      T@      `@      Z@      ,@      @     �Y@     �U@      "@      ;@     @]@      3@     �X@     �K@     �_@     �W@      @              "@      0@                      (@      @      $@      9@       @      "@      @       @      E@     �W@      @      "@     @V@      4@     �f@      1@     �d@     �B@      @              @      ?@              �?      0@      @     �D@      �?     �G@       @      @       @     �C@      P@      @       @     @R@      1@     �a@      0@     �]@     �A@               @     �O@      W@      &@      (@     �Q@      &@     �\@     �J@     �W@     �T@      @      �?      9@      :@      @      "@      @@      @     �E@      $@      K@      ?@       @      �?      9@      5@      @      @      <@      @      8@      $@      B@      9@       @                      @              @      @              3@              2@      @              �?      C@     �P@      @      @     �C@      @      R@     �E@     �D@      J@      @              0@      G@       @             �@@      @     �E@      8@      B@      A@       @      �?      6@      4@      @      @      @       @      =@      3@      @      2@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�V�GhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�n�>vW@�	           ��@       	                    �?�Ʋ �'	@           ؙ@                           �?�C+�@�           0�@                           �?�ܵ�Y�@�             l@������������������������       ��3&6VW@:            @U@������������������������       �Jΰ%O�@T            `a@                          �2@�!4�w�@�            `x@������������������������       ��C]GA@,             P@������������������������       ��Y���@�            `t@
                           �?��tF	@�           @�@                           @&�S���@�            w@������������������������       �Qzմ7�@b            `c@������������������������       �)��Y�@z            �j@                            @%B�ƹ	@�           ��@������������������������       �I�b�"�	@�            �t@������������������������       ��2)x+	@�            u@                           �?lK�	@�           ��@                           @�d�v@�           ��@                           @r��九@           �z@������������������������       ��k-K��@�            �r@������������������������       �O�4�~�	@O            �_@                           @��^*uh@�           ��@������������������������       �ю-��@�            �s@������������������������       ��:�R�]@�             t@                           @<���@�           ��@                          �2@�So#Ii@H           �@������������������������       ���B��q @�            �t@������������������������       ��(4��@~           ��@                          �8@�Dr�@�            Pp@������������������������       ���%ܒ@y            �g@������������������������       �>�#|@-            �Q@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        $@     q@     P�@      <@      J@     P|@     �X@      �@     �j@     p�@     pz@     �@@      $@     �c@      n@      5@      ?@     �n@     �K@     �m@     �a@     @o@     �m@      9@       @     �O@     �Y@      "@      @     @X@      7@     �W@      G@     @Q@     �W@      "@              9@      ;@      @      @      A@       @      K@      &@     �C@      :@                      @      &@                      *@              7@      @      6@       @                      4@      0@      @      @      5@       @      ?@       @      1@      2@               @      C@      S@      @      �?     �O@      5@      D@     �A@      >@     @Q@      "@              �?      "@                      0@      �?      *@      �?      *@      $@               @     �B@     �P@      @      �?     �G@      4@      ;@      A@      1@     �M@      "@       @     �W@      a@      (@      ;@     �b@      @@     �a@     @X@     �f@      b@      0@              8@      H@      @       @     �G@      "@     �Q@      6@     �Q@     @P@      @              *@      8@      �?              .@      @     �A@       @      F@      $@                      &@      8@       @       @      @@      @     �A@      ,@      :@     �K@      @       @     �Q@     @V@      "@      3@     �Y@      7@      R@     �R@     �[@     �S@      *@      @      ?@      @@      @      0@     �I@       @      ?@     �D@     �O@      F@      @      @     �C@     �L@       @      @      J@      .@     �D@      A@      H@     �A@       @              ]@     �s@      @      5@     �i@     �E@     ��@      R@     ��@      g@       @             �L@     �b@      @      *@     �[@      *@     0v@      8@     `o@     @T@      @              >@     �R@      �?      @      L@      $@     �Z@      ,@      V@     �C@      @              2@      L@                      B@      @      X@      @      Q@      5@                      (@      2@      �?      @      4@      @      &@      &@      4@      2@      @              ;@     @S@      @      $@     �K@      @      o@      $@     `d@      E@                      *@      <@              "@      7@      �?     �b@      @      U@      @                      ,@     �H@      @      �?      @@       @      Y@      @     �S@     �A@                     �M@     `d@       @       @     �W@      >@     y@      H@     �q@     �Y@      �?              I@     �_@      �?      @     �P@      4@     `u@      B@     `j@     �Q@                      @     �G@              �?      @       @     �d@      "@      R@      6@                      F@      T@      �?      @      N@      2@     �e@      ;@     `a@      H@                      "@      B@      �?      �?      =@      $@     �M@      (@     �Q@     �@@      �?              "@      ?@      �?      �?      0@      @     �K@      @     �G@      1@      �?                      @                      *@      @      @      @      7@      0@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�igohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?���@�	           ��@       	                    @�����@           ��@                          �8@��&ޖ@�            �@                          �3@�ۓ(�@5           �~@������������������������       ����yh@�             p@������������������������       ���J�d�@�            @m@                            �?H�t��@s            �f@������������������������       ���{�E�@<            �W@������������������������       �����`�@7            �U@
                           @�-HA�@u           ��@                          �4@6�0CO�?�            �x@������������������������       �O��U��?�            �o@������������������������       �0n�2�@Q            `a@                          �5@�$�� �@�            �i@������������������������       �aO�� @N             `@������������������������       �bS��P@3            @S@                           �?�^iv��@�           ��@                           �?X�&��	@�           (�@                          �=@o�y�"h@           y@������������������������       �l��Kb*@�            �w@������������������������       ���M��^@             9@                           �?��[Lh,
@�           ȅ@������������������������       ��<���	@�            �k@������������������������       ��M��	@0           �}@                           @�:��(�@�           �@                           �?�RY��@�            �x@������������������������       ���7�=@`            �a@������������������������       ��L��XN@�            �o@                           @��B��@�           ��@������������������������       ���K���@           x�@������������������������       �2�)G$k@�             u@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     �q@     ؀@      9@      I@     �{@     �U@     h�@     �i@     ��@     `v@     �A@       @     �S@     �c@      @      @     �[@      0@     �}@     �I@     `q@     @V@      @       @     @P@     �T@      @      @     @V@      @     `f@     �D@     �a@     �K@      @             �G@     �J@      @      @     @P@      �?      c@      6@     �Z@      @@      @              4@      6@               @      :@              U@      &@     �O@      <@                      ;@      ?@      @       @     �C@      �?     @Q@      &@     �E@      @      @       @      2@      >@               @      8@      @      :@      3@      A@      7@               @      @      2@                      @      @      @      $@      7@      4@                      &@      (@               @      3@      �?      3@      "@      &@      @                      *@     �R@                      6@      &@     pr@      $@     @a@      A@       @              "@     �H@                       @      $@     �j@      @     �U@      1@                       @      ;@                      @              c@      �?      J@      "@                      �?      6@                      @      $@     �M@       @      A@       @                      @      :@                      ,@      �?     �T@      @      J@      1@       @              @      2@                      @              M@      �?     �@@      &@       @              �?       @                      &@      �?      9@      @      3@      @              0@     @i@     �w@      6@      F@     �t@     �Q@      �@     `c@     ��@     �p@      =@      .@     @\@      d@      0@      5@     `e@     �H@     @`@     �X@     �c@     @b@      6@       @      ;@     �R@      @      @      M@      *@     @Q@      =@     �L@     �L@      @       @      9@     �R@       @      @      M@      &@     �P@      ;@      K@      G@      @               @               @                       @      @       @      @      &@              *@     �U@     �U@      (@      .@     @\@      B@     �N@     @Q@     �X@     @V@      2@      @      ;@     �@@      @              :@      *@      ,@      <@      9@      C@      "@       @     �M@     �J@      @      .@     �U@      7@     �G@     �D@     �R@     �I@      "@      �?     @V@     �k@      @      7@     `d@      5@     �{@     �L@     0x@     �^@      @              8@      Q@      �?      $@     �G@      @     �V@      B@     @R@     �C@                      @      4@      �?       @      7@       @      6@      1@      <@      2@                      1@      H@               @      8@       @      Q@      3@     �F@      5@              �?     @P@      c@      @      *@      ]@      1@     @v@      5@     �s@      U@      @      �?      D@     @[@      �?      @     �R@      $@     �q@      "@     �l@     �G@      @              9@     �E@      @      $@     �D@      @     �Q@      (@     �T@     �B@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��'hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�t�U{@�	           ��@       	                    �?X�^�!�@d           �@                          �;@��<M�@           �@                           �?�,ʁ�@�           �@������������������������       �5�4�K�@�            �j@������������������������       ���7���@:           �~@                            �?�����@Q            �^@������������������������       ��N����@+            �P@������������������������       �H�V�	@&             L@
                           �?c2r��@G           �@                            �?S�-�;@�            Pu@������������������������       �w��@A            �X@������������������������       �nG摏�@�            @n@                           �?ƥ_D�\	@u           8�@������������������������       �������@=            �\@������������������������       ��	�d�	@8           ��@                          �4@d��J#�@:           @�@                            @��G�7@C           (�@                           @ۉ���_@�           �@������������������������       ��\�!��?v           `�@������������������������       ��{_��@h            �b@                          �0@n�?�p�?e            `d@������������������������       �@`�zò�?             2@������������������������       ���@��?Z             b@                           @2��vX{@�           X�@                          �8@M��\�@@           0�@������������������������       �za�.؂@�            �u@������������������������       ���mvv@j             e@                          �?@έ؀�@�            Pr@������������������������       ���RG|@�            �q@������������������������       ��}�F��?             &@�t�b��
     h�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@     H�@      =@     �K@     �}@     �S@     ��@      h@     �@     �v@      =@      3@     `h@      s@      9@      H@      t@     �M@     �w@     @d@     �w@      o@      8@      $@     �T@     �\@      .@      *@     �^@      9@     �a@     �O@     �`@      [@      @      @     �Q@     @X@      .@      (@     @Z@      0@      a@      J@     �]@     �R@      @      �?      ,@      ?@       @      @      G@      �?     �F@      $@      E@      ,@      �?      @      L@     �P@      *@      @     �M@      .@     �V@      E@     @S@     �N@       @      @      (@      1@              �?      2@      "@      @      &@      ,@     �@@               @      @      @                      $@      @       @      $@      @      5@               @      @      &@              �?       @       @       @      �?      $@      (@              "@     @\@      h@      $@     �A@     �h@      A@      n@     �X@     �n@     �a@      5@              B@      J@              @      @@              W@      (@     �U@      9@      @              *@      1@                      "@              ,@      @     �@@      @      @              7@     �A@              @      7@             �S@      "@     �J@      2@              "@     @S@     �a@      $@      @@     �d@      A@     �b@     �U@      d@     �\@      2@      @      ,@      @              *@      <@              @      *@      9@      @      @      @     �O@     �`@      $@      3@     `a@      A@      b@     �R@      a@     @[@      ,@      �?     @U@     �j@      @      @     �c@      4@     H�@      >@     `z@     �]@      @             �A@     �X@       @      @      M@      @     `|@       @     @k@      I@      �?              >@      U@      �?      @     �G@      @     �w@       @     `d@     �G@      �?              3@     �Q@                      9@      @      u@      @     �]@      D@                      &@      ,@      �?      @      6@             �E@      @     �F@      @      �?              @      ,@      �?              &@      �?     @R@             �K@      @                                                                      .@              �?       @                      @      ,@      �?              &@      �?      M@              K@      �?              �?      I@     @]@       @      @     �X@      ,@     `l@      6@     �i@      Q@      @      �?     �D@      Q@              �?     �N@      "@     @d@      @      `@     �A@      @      �?      @@     �E@                     �F@      @     @^@       @     �R@      4@      @              "@      9@              �?      0@       @     �D@      @     �K@      .@                      "@     �H@       @      @     �B@      @     @P@      .@     �R@     �@@                      @     �H@       @      @      B@      @     @P@      ,@     �R@      <@                      @                              �?      �?              �?              @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��;EhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �3@�ݫ?r@�	           ��@       	                    �?vں���@�           ��@                           @�Ӑ�K�@           �}@                            �?���b@�            �v@������������������������       �-<R� @7            �T@������������������������       �#��t�@�            `q@                           �?��c�T�@?            �[@������������������������       �U*s�A�@            �B@������������������������       ��K�vm@*            �R@
                           �?#�ئ�@m           ��@                            �?a8İ� @1            @������������������������       �q�3�#Y@E            @]@������������������������       ���W]��@�            �w@                          �1@��o%@<           p~@������������������������       �������?�            �i@������������������������       �PA���@�            �q@                           �?�3"W�~@           4�@                           �?ɒ�|��	@�           ��@                           �?Y '�O@�            Px@������������������������       ���㞋�@J            �^@������������������������       ���jiv@�            �p@                          �;@/5'��	@�           H�@������������������������       ��RD���@d           ��@������������������������       ����D&�	@o             g@                           �?�nc��@L           ��@                            @�	�F@�            `u@������������������������       �+�&"�@�            �q@������������������������       ���黛#�?%             O@                           @���9��@j           ��@������������������������       ��_��]<@           P|@������������������������       ���>�f�@W           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     p�@      ?@     �P@     �|@      V@     �@     @k@     ��@     0v@      7@      @      V@     �i@      @      (@      `@      $@     @~@      P@     Pu@      \@      �?      @     �D@      O@      @      @     �Q@      @     �U@      D@     �W@      M@      �?      �?      7@      H@      @      @     �I@      @     @S@      5@     �S@     �G@                      �?      (@                      @              :@      @      9@      @              �?      6@      B@      @      @     �F@      @     �I@      .@      K@      D@              @      2@      ,@                      3@      �?      $@      3@      .@      &@      �?      @      (@      @                       @              @      @       @      @                      @      $@                      1@      �?      @      .@      *@      @      �?             �G@      b@      �?       @      M@      @     �x@      8@     �n@      K@                      ?@     �R@      �?      @     �D@             �g@      (@     @]@      9@                      �?      (@                      *@             �F@      @      ?@       @                      >@     �O@      �?      @      <@             @b@      @     �U@      1@                      0@     @Q@              @      1@      @     �i@      (@     @`@      =@                      @      4@                      @             �Y@      @      O@      @                      *@     �H@              @      (@      @     �Y@       @      Q@      6@              .@      l@      v@      :@      K@     �t@     �S@     �}@     @c@     �}@     `n@      6@      *@      `@      h@      3@      ?@      f@     �D@     @^@     �X@     @f@     �]@      0@              =@      L@      �?      0@      P@      @     �P@      ?@     �Q@      E@      @              5@      0@                      3@              >@      @      ;@      @       @               @      D@      �?      0@     �F@      @     �B@      <@     �E@      C@      @      *@      Y@      a@      2@      .@      \@      A@      K@     �P@      [@     @S@      $@      @     �R@     @Y@       @      "@      Y@      7@     �G@      J@     �X@      B@      @      @      :@      B@      $@      @      (@      &@      @      .@      "@     �D@      @       @      X@     �c@      @      7@     �c@     �B@     `v@      L@     �r@      _@      @              @     �D@               @     �B@      @     `a@      "@      T@      3@      @              @     �D@               @     �@@      @      Y@      @     �P@      0@      @                                              @             �C@      @      *@      @               @     @V@     �]@      @      5@     �^@      @@     `k@     �G@      k@     @Z@      @       @     �F@      K@       @       @     �P@      8@     �U@      @@     @T@     �J@                      F@      P@      @      *@      L@       @     �`@      .@      a@      J@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJM,�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��P�5;@�	           ��@       	                    �?��*G6�@^           ��@                           �?�I���@�           ܘ@                          �;@Sˋ@�@�           Ȃ@������������������������       ��h�?@S           x�@������������������������       ��	�0�|@1            �R@                           �?6��Sn	@g           ��@������������������������       �'Na��@�            `r@������������������������       ��]��	@�           ��@
                          �3@�`EOt�@s           (�@                           �?Q�n��@�            `l@������������������������       �̨ %� @2            �T@������������������������       ��h��@X             b@                          �4@ i��|@�             v@������������������������       �!i9���@)            �P@������������������������       �F�K%�@�            �q@                           �?o��מK@D           4�@                            �? YQ�!@s            �@                          �5@Ú���+�?T             a@������������������������       ���M2Q�?:            �X@������������������������       �a��Y)@            �C@                          �4@�ן�%�@           p{@������������������������       �;��1@�            `q@������������������������       ��A8f�l@n             d@                           @�����n@�           4�@                           @���<@�           @�@������������������������       ��H-�A_@-           ~@������������������������       ���\&�@�            pt@                          �<@�Rl�=@�            Pv@������������������������       ��Gx�@�            �t@������������������������       �e����S�?             6@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@     �r@     ؀@      <@     �J@     p|@     �S@     H�@     @j@     `�@     Px@      @@      *@      i@     Ps@      7@     �@@     �r@     �N@     �v@     `e@     @y@     �p@      :@      *@     �c@     @l@      2@      7@      m@      E@     @m@      `@     @r@     �h@      :@       @      E@     @V@      @      @     �U@      (@     �]@      ;@     �_@     �S@      @              B@      U@      @      @     �R@      "@     �Z@      :@      ^@      K@      @       @      @      @                      (@      @      *@      �?      @      9@              &@      ]@      a@      ,@      0@     @b@      >@     �\@     �Y@     �d@     �]@      3@              3@      I@      �?      @      A@      �?     �I@      >@     �P@     �A@      �?      &@     @X@     �U@      *@      &@      \@      =@      P@      R@     �X@      U@      2@              E@     �T@      @      $@     @Q@      3@     �_@      E@      \@      R@                      0@      B@                      3@             �L@      0@     �M@      8@                      $@      @                      @              4@      �?      C@      @                      @     �@@                      *@             �B@      .@      5@      4@                      :@     �G@      @      $@      I@      3@     �Q@      :@     �J@      H@                              $@      @      @      .@      @      &@       @      @      $@                      :@     �B@              @     �A@      ,@     �M@      8@      H@      C@                     �Y@     �l@      @      4@     @c@      1@      �@     �C@     �y@     �]@      @              4@     �S@              @      <@      @     �q@      @     �_@      6@      �?                      (@                      @       @     @T@              ?@      @                              @                      @              P@              8@      @                               @                      @       @      1@              @      �?                      4@     �P@              @      5@      @     @i@      @      X@      2@      �?              .@      D@              @       @             @a@      @      M@       @      �?              @      ;@                      *@      @      P@      �?      C@      $@                     �T@     �b@      @      .@     �_@      (@     Pv@     �@@     �q@     @X@      @             �L@     �\@              @      V@      @     @q@      2@     �g@     �K@      @              C@     �P@               @     @P@      @     �a@      .@      Z@      E@      @              3@      H@               @      7@             �`@      @      U@      *@                      :@      B@      @      &@      C@       @     @T@      .@     @W@      E@       @              3@      B@      @      &@     �A@       @     @T@      .@     @V@      A@       @              @                              @                              @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��1hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @3�� �N@�	           ��@       	                    �?��E~H�@x           <�@                           �?��3�-	@           l�@                          �6@�d:4@;           �~@������������������������       �љ���@�            �r@������������������������       ��UΜ_�@v            @g@                           �?�V�^�	@�           ̑@������������������������       ��`+5��	@�            `w@������������������������       �	���K	@�           �@
                            @��
@l           �@                            �?!�I�@           �y@������������������������       �-g8r�@t             h@������������������������       ���M#w�@�            �k@                          �5@��`��3@e            �d@������������������������       �@���c@6             V@������������������������       �����@/            �S@                           �?:d ^@8           ��@                          �5@?��E�� @x           X�@                           @J��*�v�?           `y@������������������������       �& L�v#@=             W@������������������������       ����˘�?�            �s@                           �?�H��Y@s            �f@������������������������       �e�?d@B            �Y@������������������������       ���Z$3@1            �S@                           @=)#p5K@�           ��@                          �1@��O��@�           �@������������������������       ��Zi6�y�?~            @i@������������������������       ��2�P�@,           ��@                           @��W}Z@             ?@������������������������       ��swn`P@
             .@������������������������       �>��_�@             0@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     �r@     x�@      B@      J@     `|@     �T@     ��@     �j@     ��@     0w@     �@@      $@     �i@     �s@      9@     �B@     �s@     �O@      w@     `f@     �w@      q@      ?@      $@     �d@      n@      9@      ?@      o@      I@     �m@     �^@     pp@     �i@      <@              L@     �R@      @      @     �K@      @     @[@      =@     �W@     �I@      @              D@     �C@       @      �?      8@       @     @W@      4@      M@      5@       @              0@      B@       @      @      ?@      �?      0@      "@     �B@      >@       @      $@     @[@     �d@      5@      8@      h@     �G@      `@     �W@      e@     `c@      8@      @      @@     �Q@      &@      @     �Q@      6@      A@      9@      A@     �J@      .@      @     @S@      X@      $@      4@     �^@      9@     �W@     @Q@     �`@     �Y@      "@             �C@      S@              @      Q@      *@     �`@      L@     �]@     �P@      @              7@     �G@              @      K@      (@     @V@      F@     �W@     �E@      @              @      <@              @      5@      @     �I@      ,@     �D@      6@      @              1@      3@              �?     �@@       @      C@      >@     �J@      5@                      0@      =@               @      ,@      �?      F@      (@      9@      7@                       @      4@               @      @      �?      @@      @      &@      "@                      ,@      "@                      "@              (@      @      ,@      ,@               @     �W@     @n@      &@      .@     @a@      3@     ��@      B@     �y@     �X@       @              0@     �U@              �?     �D@      @     Pq@      @     �`@      6@                      (@      N@              �?      5@             �k@      @     @S@      "@                       @      3@                      @              D@              1@      @                      @     �D@              �?      1@             �f@      @      N@      @                      @      ;@                      4@      @      K@      @      L@      *@                      @      .@                      @      �?     �C@      �?      =@      @                      �?      (@                      *@       @      .@      @      ;@      @               @     �S@     `c@      &@      ,@     @X@      0@     �v@      =@     @q@     @S@       @       @     @R@      c@       @      *@     @V@      *@     pv@      <@     0q@     �R@       @              @      9@              �?      "@             @Z@      @      H@      @               @     �Q@      `@       @      (@      T@      *@     �o@      7@     `l@      Q@       @              @       @      @      �?       @      @      @      �?      �?      @                       @              @              @       @              �?              �?                      @       @              �?       @      �?      @              �?       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJo�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�9��_|@�	           ��@       	                   �2@��@X�	@o           r�@                           �?�-~���@,           �}@                            �?�m�j�g@n            �d@������������������������       ��ŁaV�@!             K@������������������������       �9F'�m@M            �[@                            @5
uC�@�            `s@������������������������       ��8خ�@s            �f@������������������������       ��|�&�@K             `@
                           �?s��X!v	@C           |�@                            �?�ҟ~W�@,           �|@������������������������       ������@�            pp@������������������������       ���PI��@�            @h@                           �?�Y�{��	@           X�@������������������������       �a�YВ<
@W           ��@������������������������       �*��K>�@�             t@                          �4@��F�@           @�@                           �?�5o�@7            �@                          �3@s�a�B��?�            Pw@������������������������       ��^&i��?�             s@������������������������       �M��`�w @*            @Q@                           @�_1��@T           x�@������������������������       ��cY��@0           @������������������������       ���!j�@$             O@                          �8@S9S@�           `�@                          �5@[\e�a@#           �{@������������������������       ����t�@\            �a@������������������������       �����@C@�             s@                          �:@d9�j��@�            �r@������������������������       �(78��L@N             `@������������������������       ��% [I�@o            �e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     �q@     X�@      B@     �I@     �z@     �V@     x�@      l@     H�@     Py@      B@      3@     `i@     @v@     �@@     �A@      r@     �P@     x@     �g@     �u@     pq@      >@       @      3@     �Q@      �?      @      G@      @     `c@      D@     @U@     �F@       @       @      @      :@      �?              7@      �?      L@      (@      8@      ,@      �?                      1@                      @              1@      @      &@      �?      �?       @      @      "@      �?              4@      �?     �C@       @      *@      *@                      .@     �F@              @      7@      @     �X@      <@     �N@      ?@      �?              @      7@                      (@      @     �M@      6@     �C@      0@      �?              "@      6@              @      &@      �?      D@      @      6@      .@              1@      g@     �q@      @@      @@     �n@     �N@     �l@     �b@     `p@     @m@      <@              G@      R@       @      @     �K@       @     �W@      5@     @Y@     �I@      @              <@      F@      �?      @      7@              J@      "@     �P@      =@      @              2@      <@      �?       @      @@       @     �E@      (@      A@      6@              1@     @a@     �j@      >@      9@     �g@     �M@     �`@      `@      d@     �f@      7@      1@     �Z@     �b@      =@      1@     �a@     �I@     �V@     �X@     �Z@     �b@      7@              @@      O@      �?       @     �G@       @      F@      >@      K@      A@              �?      T@     �h@      @      0@     @a@      8@     p�@     �A@     �z@     �_@      @              D@     @V@       @       @      J@      @     �z@      "@      n@      K@       @              $@      ?@              @      2@             �j@      @     @T@      &@       @              "@      6@               @      &@             �e@      @      R@      @       @              �?      "@               @      @             �B@              "@      @                      >@      M@       @      @      A@      @     @k@      @     �c@     �E@                      :@      H@       @      @     �@@      @     @h@      @     �b@     �@@                      @      $@                      �?              8@       @      &@      $@              �?      D@     �[@      �?       @     �U@      2@      h@      :@     �g@      R@      @      �?      7@     �T@      �?      @      H@      .@      `@      @     �Z@      <@      @               @      ;@               @      ,@       @     �A@      �?      F@      @      @      �?      5@     �K@      �?      �?      A@      @     �W@      @     �O@      5@      �?              1@      <@              @      C@      @     �O@      4@     �T@      F@                       @      @                      *@       @      ?@      @      F@      8@                      .@      5@              @      9@      �?      @@      .@     �C@      4@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�q��7�@�	           ��@       	                    �?@޶�>�	@           ��@                           �?:��@�           ��@                          �:@�i�@��@�             o@������������������������       ����\�@�            @i@������������������������       �~�/%�@            �G@                            �?&4
��@�            `v@������������������������       �����@�            `n@������������������������       ��kb��w@K            �\@
                           �?~zv�	@�           4�@                           �?Ӻi|1
@�            �u@������������������������       �k~hPm	@^            `a@������������������������       �f�Rr�	@�            `j@                          �<@�4٬Z�	@�           x�@������������������������       ���B�7	@k           h�@������������������������       ����Tt	@B            �X@                           �?TMZ���@�           ��@                            �?ں3��@�           �@                          �8@�f��uO @|             g@������������������������       ��\����?n            @d@������������������������       �z��-@             6@                          �8@�����@f           H�@������������������������       ��n��@3           �@������������������������       ���J���@3            �S@                          �1@&
̨�@�           p�@                           @�@7��@�            0p@������������������������       �_z��K�@'             M@������������������������       ��U㑑� @�             i@                            �?�/�+�@           d�@������������������������       ����R�@�           @�@������������������������       �^K�'�N@T           ��@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        5@     �s@     Ȁ@      B@      P@     �{@      V@     0�@      j@     (�@      v@      D@      5@     �g@     �o@      8@      E@     p@     �H@     `i@     �_@     �o@      h@      ?@      @      G@     �Z@      @      .@     �V@      "@     �\@     �E@     �Y@     �P@      @      @      3@     �H@       @      @     �E@       @      J@      *@      ?@      :@       @      @      0@      C@       @      @      @@       @      J@      "@      <@      *@       @       @      @      &@                      &@                      @      @      *@                      ;@      M@       @      $@      H@      @      O@      >@      R@      D@       @              2@     �B@       @      @      ;@      @     �E@      1@      J@     �A@      �?              "@      5@              @      5@       @      3@      *@      4@      @      �?      0@      b@     @b@      4@      ;@     �d@      D@     @V@     �T@      c@     �_@      ;@      @     �J@     �G@      &@      $@     �I@      1@     �B@     �@@     �@@      H@      @              0@      ,@       @      @      2@      @      ;@      ,@      *@      4@       @      @     �B@     �@@      "@      @     �@@      &@      $@      3@      4@      <@      @      (@      W@     �X@      "@      1@     �\@      7@      J@      I@     �]@     �S@      5@      (@      U@     �V@      @       @     �X@      4@      H@      B@     �[@     �L@      0@               @       @       @      "@      0@      @      @      ,@       @      5@      @             �^@     �q@      (@      6@     `g@     �C@     �@     �T@     0�@      d@      "@              ?@      U@              @     �@@      &@     �w@      ,@     �d@      C@      @              �?      1@               @      @      @     @Y@             �B@      $@      @              �?      0@               @      @      �?     �W@             �A@      @                              �?                              @      @               @      @      @              >@     �P@               @      :@      @     �q@      ,@     @`@      <@      �?              >@      N@               @      6@       @      p@      &@     �Y@      2@      �?                      @                      @      @      7@      @      <@      $@                     �V@      i@      (@      2@     @c@      <@     0|@     @Q@     �u@     �^@      @              @     �E@               @      @             @Z@      "@     �Q@      1@                       @      *@                       @              2@      @      (@      @                      @      >@               @      @             �U@      @     �M@      (@                     @U@     �c@      (@      0@     �b@      <@     �u@      N@     �q@     @Z@      @             �M@      T@      @      @     �R@      0@      f@      B@     `d@     �O@       @              :@     @S@      "@      "@     @R@      (@     @e@      8@     @]@      E@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?Q�A��E@�	           ��@       	                    �?8��ؐ@           |�@                          �7@��I��@2           0~@                           �?����8@@�             s@������������������������       ��7��� @L            @_@������������������������       ��MK,�@{            `f@                           �?u��k��@k            `f@������������������������       ��g�n�S@3             U@������������������������       ����Ű@8            �W@
                          �>@	�Lv��@�           ��@                           @�m�H&@�           H�@������������������������       ��I��א@Y           �@������������������������       �����@~             i@������������������������       �����|'@             3@                          �5@����.@�           Ԥ@                            �?mk���@e           ؕ@                          �4@y��!�@�            �t@������������������������       �z��;��@�            �q@������������������������       �H`��>@%             K@                          �1@���g@�           ��@������������������������       �?�3��%@�            `r@������������������������       �����@�           �@                           @��Be	@"           Г@                            �?�Ϙ�˖	@           ��@������������������������       �PX��!
@           �y@������������������������       ���v荑@�            �y@                           @0�ܡl�@           �{@������������������������       ��J
��@�            �p@������������������������       �ڊ���n@v            @f@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        3@      t@     ��@      8@      G@     p}@     �S@     �@     �j@     X�@     �w@     �A@       @      U@     �d@      @      @      ^@      $@     p|@     �C@      q@     �T@      @       @      I@      Q@      �?      @     �O@       @     �_@      7@     �V@      G@      @              A@     �B@              �?      ;@       @     �W@      *@     �Q@      6@      @              "@      *@                      @              J@       @     �C@      @                      9@      8@              �?      4@       @      E@      &@      @@      3@      @       @      0@      ?@      �?      @      B@             �@@      $@      3@      8@      �?       @      "@      .@      �?      @      *@              "@      @      "@      0@                      @      0@              �?      7@              8@      @      $@       @      �?              A@     �X@       @             �L@       @     �t@      0@     �f@      B@       @              @@     �X@       @              J@       @     `t@      &@     �f@      @@       @              <@      O@                      A@       @     �o@      @     @`@      9@      �?              @     �B@       @              2@             @R@      @     �I@      @      �?               @                              @               @      @      �?      @              1@     �m@     �v@      5@     �C@     �u@     @Q@     ��@     �e@     �@     `r@      =@       @     @T@     `i@      "@      1@     @e@      <@     @w@     @R@     �r@     �^@      &@              2@      E@               @     �A@      @     @Z@      ,@     �R@      ?@       @              .@      =@              �?     �A@      @     @V@      ,@     �M@      <@       @              @      *@              �?               @      0@              0@      @               @     �O@      d@      "@      .@     �`@      7@     �p@     �M@     �l@      W@      @      �?      0@      F@      �?      �?      :@             @X@      *@      S@      3@              @     �G@     @]@       @      ,@     @[@      7@     @e@      G@      c@     @R@      @      "@     `c@     �c@      (@      6@     �f@     �D@     @h@     �Y@     �i@     `e@      2@      "@     @]@     @Y@      $@      ,@      `@     �A@      V@     @T@      X@     �_@      1@      @     �J@     �H@      @      *@     �K@      7@      D@     �K@     �F@     �M@      @       @      P@      J@      @      �?     �R@      (@      H@      :@     �I@     �P@      &@              C@      M@       @       @      J@      @     �Z@      5@      [@     �F@      �?              .@      @@               @      6@      @     �Q@      (@     �R@      ;@                      7@      :@       @              >@             �A@      "@      A@      2@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJkwdhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�� �|s@�	           ��@       	                   �1@���@[           �@                          �0@��!�R@�           ��@                            @��$��@w            �f@������������������������       �-�O��� @a             c@������������������������       ���dN@             >@                           @� �[��@           �{@������������������������       �l 0���@�            �s@������������������������       ����Ԥ_@P             _@
                           @�{�CC@�           �@                           �?Q�o��@           ��@������������������������       ����ϐ�@�            �r@������������������������       ��9���u@T           �@                           @��w��3@�           x�@������������������������       ��Mn���@V           p�@������������������������       �<�E�ߙ@e             d@                           �?�/u��@G           \�@                          �=@_p��O@#           �|@                          �7@�����@	           0z@������������������������       �-h�wi2@W            �`@������������������������       �g��M�*@�            �q@                            @�몚�~@             D@������������������������       ����D3l@             5@������������������������       ���'�,�@
             3@                           @'G�L	@$           0�@                          �6@�4�{�	@           ��@������������������������       ��<��@[            �c@������������������������       �M�Y���	@�           ��@                           @���r�@           �{@������������������������       �vy�@f@           �z@������������������������       ��O�kS@             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        *@      t@     X�@      @@      M@      {@     �T@     x�@     �m@     ��@     px@      ;@      @      _@     @r@      ,@      3@     �i@      :@      �@     �W@     `~@     �f@      "@       @      9@      T@       @      @      C@      �?     pp@      6@     �a@     �E@       @              @      >@              �?      ,@             �U@      @      >@      ,@                      @      <@                      &@              R@              :@      (@                      �?       @              �?      @              ,@      @      @       @               @      5@      I@       @      @      8@      �?      f@      3@     �[@      =@       @       @      0@     �D@       @              2@      �?     �_@      .@     @Q@      =@                      @      "@              @      @             �I@      @      E@               @      @     �X@     �j@      (@      *@      e@      9@     �{@      R@     �u@     `a@      @      @     �Q@     �]@      $@      @     @_@      3@     �e@      P@     `d@     �W@       @      �?      ;@     �K@      @       @     �E@      $@     �Q@      ;@      F@      3@               @      F@     �O@      @      @     �T@      "@      Z@     �B@     �]@     �R@       @              <@     �W@       @      @      F@      @     �p@       @     �f@     �F@      @              (@     �R@      �?      @      A@       @      l@      @      a@      >@                      0@      3@      �?              $@      @     �E@       @      G@      .@      @       @     �h@     pp@      2@     �C@     `l@      L@     �p@      b@     �r@      j@      2@      �?      F@     �S@      �?      "@     �G@      @      X@      9@     �X@     �G@      @      �?     �E@     �R@      �?      @     �D@      @     �W@      *@     �W@     �D@      @              .@      8@      �?              (@             �C@              6@      3@              �?      <@     �I@              @      =@      @     �K@      *@      R@      6@      @              �?      @              @      @      �?       @      (@      @      @                      �?       @                      @      �?              @      @      @                               @              @      @               @      @       @      �?              @     @c@      g@      1@      >@     �f@     �H@     �e@      ^@      i@     @d@      ,@      @     �]@     @`@      &@      :@     �^@      G@     @R@     �W@      [@     �X@      ,@      @     �@@      5@      �?      "@      3@      @      1@      5@      4@       @              @     �U@     @[@      $@      1@     �Y@     �E@      L@     @R@      V@     �V@      ,@             �A@      K@      @      @      M@      @     �Y@      :@      W@     �O@                      <@      J@      @      @     �K@      @     �Y@      6@     �V@     �O@                      @       @      �?              @                      @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @��I#�@�	           ��@       	                   �5@�6m���@�           ��@                           �?rR�L@�           �@                          �1@�D��@�           ��@������������������������       ���G�]T@x             j@������������������������       ��)��=	@�           0�@                            �?��g��@�             t@������������������������       �j����@;            �V@������������������������       ��@�Ǽ@�             m@
                           @�Bv'	@�           4�@                           �?��t���@r           H�@������������������������       �*f��f�@�             t@������������������������       �$��;&U	@�           8�@                           @XV���@A             Y@������������������������       ���ھ�b@.            �Q@������������������������       �Bإq�6@             =@                           @�j��@/           �@                            �?��@�           ��@                          �1@Im3�@�           ��@������������������������       �V�rF1d�?b            `d@������������������������       �V}Rqu�@%           P}@                            @���3�@U           `@������������������������       �'Y���@�            v@������������������������       �3��#� @a            �b@                           �?���S�@S           ��@                            @����@�            �p@������������������������       �'���&�@z             h@������������������������       �3�����@2            @S@                            �?���t��@�            �p@������������������������       �S��}�@'             N@������������������������       �����@�            �i@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �t@      �@      B@     �K@     �~@     �R@     ��@      l@     ��@     �v@      >@      4@     �o@     �r@      =@     �C@     �v@      M@     @u@     �g@     �w@     p@      :@       @     �V@     @a@      *@      4@     @d@      ;@     @m@     �V@      m@     �]@      &@       @     @R@     �V@       @      .@      _@      5@     �b@     @Q@     �c@     �W@      &@              *@      6@       @      @     �@@      �?     �H@      $@      H@      ;@               @      N@     @Q@      @      &@     �V@      4@     @Y@     �M@     �[@      Q@      &@              1@     �G@      @      @      C@      @      U@      6@     �R@      8@                      @      &@              �?      @      @      :@      @      9@      (@                      *@      B@      @      @     �@@      @      M@      3@     �H@      (@              (@     @d@      d@      0@      3@     �h@      ?@     �Z@     �X@      b@     @a@      .@      "@     @b@     �b@      0@      3@     �f@      :@     �X@     @S@     �`@     �`@      &@       @     �H@      H@       @      @      L@       @      E@      0@     �L@      D@      @      @     @X@     �Y@      ,@      .@     @_@      8@     �L@     �N@     �S@      W@      @      @      0@      &@                      1@      @      @      5@      $@      @      @       @      (@      &@                      (@      @      @      *@       @      @      @      �?      @                              @      �?               @       @      �?      �?       @     @T@      k@      @      0@     �`@      1@     �@      B@     py@      [@      @       @     �K@      a@      �?      @     �S@      (@     `~@      1@      q@     @P@       @              ;@     �V@      �?       @     �@@      @     pp@      &@     @c@      F@      �?              @      *@                      @             �Z@              <@      @                      7@     �S@      �?       @      ;@      @     �c@      &@     �_@     �C@      �?       @      <@      G@              @     �F@      @     �k@      @      ^@      5@      �?       @      7@     �B@              @      C@      @     �c@      @     �Q@      0@      �?              @      "@                      @      @     �P@      @      I@      @                      :@      T@      @      &@     �L@      @     �b@      3@     �`@     �E@       @              (@      D@      @      $@      >@      �?     �S@      @     @P@      6@                      &@      ?@      @      @      :@              H@      @     �H@      (@                      �?      "@              @      @      �?      ?@       @      0@      $@                      ,@      D@      @      �?      ;@      @      R@      (@      Q@      5@       @              @      @      �?              @       @      9@      @      *@      @                       @     �B@       @      �?      8@       @     �G@      "@     �K@      1@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJmp5{hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@\��� @�	           ��@       	                    �?�K�ă@V           Ơ@                           @	"����@�            �@                          �4@m)=KT@i           8�@������������������������       ��h&�%�@*            ~@������������������������       �|���@?            @Y@                           @�n�ް@	@k            �c@������������������������       �%,���	@L            �Z@������������������������       �E��r��@            �I@
                           @�Cȷs@�           ��@                          �1@�nR�@t           ��@������������������������       �$IT��B @o             f@������������������������       ���IN�@           0z@                           �?l,Vt�'@           `�@������������������������       ��]-�0��?�            �q@������������������������       �|���@V           ��@                           �?:��?${@Y           ��@                          �:@<N�	@-           ��@                           @"���72	@c           ��@������������������������       �-Zeg	R@�            �u@������������������������       �7+�o.�	@�             k@                          �?@<�Ϥ�@	@�            pt@������������������������       ���Ev6	@�            @o@������������������������       ��o�;@*            @S@                          �8@g�_!�@,           8�@                           @����@           `z@������������������������       ���<CN�@L            �^@������������������������       ��2>x�h@�            �r@                           @��	�ޕ@           |@������������������������       ���
�1@           �z@������������������������       �Q�V#k@
             2@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     @r@     �@      4@     �N@      {@     @S@     ��@     �m@      �@      u@      :@      @     @^@     `q@       @      @@     �h@      @@     Ȇ@     @X@     @~@     �b@      $@      @     �O@      W@      @      0@     �Z@      &@     @a@     �H@     @e@      S@       @      @      F@     �P@      @      (@     @R@      @     �^@      ?@      c@     @P@       @      @     �E@      I@      @      @      P@      @     �[@      8@      ^@     �J@       @      �?      �?      0@      �?       @      "@      �?      *@      @      @@      (@               @      3@      :@      �?      @     �@@      @      .@      2@      2@      &@      @              ,@      1@      �?      @      2@       @      (@      .@      (@       @      @       @      @      "@                      .@       @      @      @      @      @      @              M@     @g@      @      0@     @W@      5@     x�@      H@     �s@     �R@       @              ?@      Y@              @     �D@      1@     @l@     �@@     @[@      >@      �?              @      2@                       @             �X@       @      :@      &@                      9@     �T@              @     �@@      1@     �_@      9@     �T@      3@      �?              ;@     �U@      @      "@      J@      @     �v@      .@     �i@     �F@      �?              @     �@@               @       @             @e@      @      M@      @                      7@     �J@      @      @      F@      @     `h@      &@     `b@     �D@      �?      0@     `e@     �p@      (@      =@     `m@     �F@     �t@     �a@     �s@      g@      0@      .@     �[@     �`@      $@      3@     �`@      ?@     �Y@     @U@     �`@     @[@      *@       @     �R@      X@      @      .@     @T@      4@     @R@     �K@     �V@     �E@      $@              F@      I@      @       @      M@      &@      J@      9@     �Q@      :@      @       @      ?@      G@      @      @      7@      "@      5@      >@      5@      1@      @      *@      B@      B@      @      @     �J@      &@      >@      >@      E@     �P@      @       @      3@      >@      �?      @     �C@      &@      ;@      7@      A@     �I@      @      @      1@      @       @              ,@              @      @       @      .@              �?      N@      a@       @      $@     @Y@      ,@     �l@      L@     �f@      S@      @      �?      A@     �R@       @      @     �J@       @      ]@      ,@      T@     �C@       @              *@      6@               @      3@              8@      @      3@      1@      �?      �?      5@     �J@       @       @      A@       @      W@       @     �N@      6@      �?              :@      O@              @      H@      (@      \@      E@     �Y@     �B@      �?              7@     �N@              @     �E@      @      \@      E@      Y@     �B@      �?              @      �?                      @      @                      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ� ehG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�)�.O@�	           ��@       	                    �?�BIͦ�@�           d�@                          �5@膄�#	@           ��@                          �0@�ѐ�<@�           ��@������������������������       ��jm1�~@!             K@������������������������       �����O@�           �@                          �;@W�/�	@2           x�@������������������������       �Tϣ0�@�           ��@������������������������       ��H��!
@�            �o@
                           �?
��W�D@~           ��@                          �;@	�<��@q             e@������������������������       ��:��=x@h            `c@������������������������       �Nɱ���@	             ,@                          �3@)?Oӥ@           pz@������������������������       �S|6W�@Y            `a@������������������������       ����y@�            �q@                           @X��ֆ@#           \�@                           �?�*�-��@           ��@                          �4@+Xx�o@g           ��@������������������������       �	��oI��?�            pu@������������������������       �C�@�            �k@                          �7@�k����@�           $�@������������������������       �kR�U@�           X�@������������������������       �#�:W�@�            �q@                            �?l</?
�@             8@������������������������       �+�%W�@	             0@������������������������       �       @              @�t�bh�h5h8K ��h:��R�(KKKK��h��B 
        1@     r@     H�@      <@     �J@     }@      T@     ��@     �l@     �@      v@     �B@      .@     �j@     �u@      5@     �B@     �s@      O@     0w@     �f@     �w@      n@     �@@      .@     @d@     `p@      4@      =@     �m@     �G@      l@     @a@      q@     �h@      ;@       @      L@     �\@      $@      $@     �[@      3@     �`@      H@     �c@     �T@      @              �?      ,@               @      3@              @      �?      @      @               @     �K@      Y@      $@       @     �V@      3@     �_@     �G@      c@     �S@      @      @     �Z@     �b@      $@      3@      `@      <@     �V@     �V@      ]@     �\@      6@             �Q@      ]@      @      *@     �X@      1@     �R@      P@     �U@      P@      ,@      @     �A@      @@      @      @      =@      &@      0@      :@      =@     �I@       @             �J@      V@      �?       @     �S@      .@     `b@     �F@     @[@      E@      @              .@      .@                      0@      �?      O@      @     �H@       @      @              (@      *@                      ,@      �?     �N@      @     �H@      �?                      @       @                       @              �?       @              �?      @              C@     @R@      �?       @      O@      ,@     @U@     �C@      N@      D@      @              "@      .@              �?      0@      @      H@      (@      7@      (@                      =@      M@      �?      @      G@      &@     �B@      ;@     �B@      <@      @       @     �R@     `i@      @      0@     �b@      2@     ��@     �F@     0z@      \@      @       @     �Q@     `i@      @      *@      b@      *@     ��@      E@      z@      \@      @              (@     �Q@      �?      �?      @@      @     �p@      .@      a@      ;@      �?              @      ?@              �?      "@              h@      @     �T@      .@      �?              @     �C@      �?              7@      @     @R@      "@     �K@      (@               @     �M@     �`@      @      (@      \@      "@      w@      ;@     �q@     @U@      @             �B@     �Y@      @       @      P@      @     �s@      *@      j@      I@      @       @      6@      ?@      �?      @      H@      @     �J@      ,@      R@     �A@                      @               @      @      @      @       @      @      �?                               @               @      @      �?      @      �?       @                                      �?                              @              �?      �?      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJi
uhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �6@z(�c@�	           ��@       	                    �?�?I��-@           D�@                           @ްȐ$=@�           l�@                            �?��~�@�@-           }@������������������������       �/�a�7	@�             o@������������������������       ���!�K@�             k@                           �?>�l��E@�           P�@������������������������       ��
2@�" @�             o@������������������������       ���}��@�             y@
                           �?H�O�@S           �@                            �?{}o��A@�            x@������������������������       ��%�x�= @K            �]@������������������������       ��=]�� @�            �p@                          �1@k�5��@\           0�@������������������������       ���r��@u            `i@������������������������       ��RWb@�           ؇@                          �;@�U�EҦ@�           ��@                           �?�	t:@�           �@                            �?ۥr�	@1           0}@������������������������       �?.��P1@p            @e@������������������������       ���%��<	@�            �r@                          �9@��*�Tc@[           ��@������������������������       �>%�z̓@�            �v@������������������������       �EQ`n�D@w            `h@                           �?G*[��@           @z@                          �?@��$�	@�            0p@������������������������       �⬛!i@|             i@������������������������       ��(�7�!	@'            �M@                           �?���SC@k             d@������������������������       � �aQ��@.            �R@������������������������       ���r��@=            �U@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     �@      @@      I@     �}@      U@     ��@     @m@     0�@     �u@      :@      *@     �b@     �u@      ,@      =@     pp@      J@     �@     @]@     `�@     �f@       @       @     �Q@     �a@      "@      .@     @`@      ;@     �w@     �H@     �i@     �R@      @       @     �D@     @S@       @      $@     @Q@      2@     �V@     �@@      R@      D@      @      @      6@      H@              "@      B@      @     �A@      8@     �A@      7@      @       @      3@      =@       @      �?     �@@      &@      L@      "@     �B@      1@                      >@     �O@      @      @     �N@      "@      r@      0@     �`@     �A@                      @      :@               @      3@      @      b@      @     �A@       @                      8@     �B@      @      @      E@      @     @b@      (@     �X@      ;@              @     �S@     �i@      @      ,@     �`@      9@     Px@      Q@     �s@     @Z@      @              8@     @P@              �?      @@             `a@      "@     @W@      5@      �?              @      9@                      @              H@             �@@      @                      2@      D@              �?      =@             �V@      "@      N@      1@      �?      @      K@     �a@      @      *@     @Y@      9@     @o@     �M@      l@      U@      @              (@      =@                      .@             �P@      "@     �J@      2@              @      E@     @\@      @      *@     �U@      9@     �f@      I@     �e@     �P@      @      "@     @c@     �h@      2@      5@      k@      @@     �j@     @]@     �q@      e@      2@      @     �Y@     `b@      ,@      .@     �a@      1@     `f@      T@      k@      X@      ,@      �?     �N@      R@      *@      "@     @W@      $@      H@     �F@     @Q@      A@      (@              =@      8@       @      @     �@@      @      4@      6@      3@      *@      �?      �?      @@      H@      &@      @      N@      @      <@      7@      I@      5@      &@       @     �D@     �R@      �?      @      I@      @     ``@     �A@     �b@      O@       @       @      9@     �K@              @      E@      @      V@      .@     @U@     �D@       @              0@      4@      �?       @       @      �?     �E@      4@     �O@      5@              @      J@      J@      @      @     @R@      .@     �@@     �B@     @P@     @R@      @      @      @@      9@      @      @     �C@      (@      .@      :@      @@     �N@       @      @      3@      3@      @      �?      >@       @      .@      7@      ;@     �I@               @      *@      @      �?      @      "@      @              @      @      $@       @              4@      ;@              �?      A@      @      2@      &@     �@@      (@       @              $@      ,@              �?      .@      �?      (@      @      .@      �?                      $@      *@                      3@       @      @      @      2@      &@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ\�<thG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@ں2.V@�	           ��@       	                     �?]�����@|           ,�@                           @�x�<�H@k           8�@                          �1@>	T�@           x@������������������������       �Z�����@E            @[@������������������������       ���fG^d@�            @q@                           @��<��?g            �d@������������������������       �p	��r�?%            �K@������������������������       ��]ؠ� @B            �[@
                          �1@����'@           ��@                           @�b�;��@           `{@������������������������       �-|d�� @�            �l@������������������������       ���rm�@�             j@                           @k��7@�           �@������������������������       �Vi�X-@�           Ї@������������������������       ����â@           �{@                          �<@��nP��@G           ̚@                           �?�g�PT@q           ��@                           �?�b`O�	@�           ��@������������������������       ��=���@�            �n@������������������������       �iU��;/
@	           �y@                           @$f;@�           ��@������������������������       �r��p*@�            �j@������������������������       ��=\\?@B           �@                           �?Ia�{	@�            0u@                          �>@3A�5Z�@:            �W@������������������������       ���u��@             F@������������������������       �w���i"@             I@                            @hv��qh	@�            �n@������������������������       �Z\�V�1@c            `c@������������������������       �0Q�X��	@9            �V@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     Ѐ@      6@     �P@     �|@     @U@     ��@     �k@     @�@     0v@      ?@      $@     @a@      r@       @      5@     �m@      @@     ��@     @V@     �|@     �e@      *@              ?@      L@              �?     @P@      @      i@      9@      `@     �B@      @              =@     �H@              �?      F@      @     �\@      8@     @U@      ?@      @               @      *@                       @              I@      @      0@       @                      5@      B@              �?      B@      @      P@      2@     @Q@      7@      @               @      @                      5@             �U@      �?     �E@      @                                                       @             �C@              ,@                               @      @                      3@             �G@      �?      =@      @              $@     �Z@     @m@       @      4@     `e@      ;@     h�@      P@     �t@      a@      $@              ;@     �I@                     �A@             `g@      2@      X@      6@       @              *@      .@                      1@             @_@      &@      C@       @       @              ,@      B@                      2@              O@      @      M@      ,@              $@      T@     �f@       @      4@      a@      ;@      u@      G@     �m@     �\@       @      $@     �N@     �_@       @      0@     �Z@      :@     �c@     �B@     �a@      R@      @              3@     �L@      @      @      =@      �?     �f@      "@     �X@      E@      �?      "@     @f@      o@      ,@     �F@     �k@     �J@     �t@     �`@     �q@     �f@      2@      @     �b@     �h@       @      >@     @e@     �B@     �r@     �X@     �m@     �^@      0@      @     �V@     �X@      @      6@      Z@      4@     �U@     �P@      T@      O@      ,@      �?      @@     �E@              @      G@      @      F@      (@      C@      2@      @      @     �M@     �K@      @      0@      M@      1@      E@     �K@      E@      F@      $@             �M@     �X@      @       @     �P@      1@      k@      @@     �c@      N@       @              ?@      >@               @      ;@       @     �H@      $@      D@      .@       @              <@     @Q@      @      @     �C@      "@     �d@      6@     �]@     �F@               @      <@     �I@      @      .@     �I@      0@      ?@      A@     �E@      N@       @              @      0@               @      &@      �?      $@      "@      ,@      4@       @               @      (@               @                      @      �?       @      &@       @              �?      @              @      &@      �?      @       @      @      "@               @      9@     �A@      @      @      D@      .@      5@      9@      =@      D@                      .@      2@      @       @      @@      *@      $@      ,@      0@      @@               @      $@      1@      @      @       @       @      &@      &@      *@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��-hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��~�S@�	           ��@       	                    �?[�lY=@           0�@                           �?�)J>�q@7           p~@                          �5@z�]d�@u            �g@������������������������       �t��-�N@E             [@������������������������       ���g��@0             T@                           �?p�,hV@�            �r@������������������������       ����_�@`             c@������������������������       �٨բi�@b            @b@
                            �?n<���@�           (�@                          �9@qJ��?� @y            `h@������������������������       ����m� �?p            @f@������������������������       ��߇�@	             1@                           >@x�Gg=�@]           �@������������������������       �n���n@T           ��@������������������������       ���h%vO@	             ,@                           @$���L@�           ��@                           @K�F��w	@�           ��@                          �3@w@��PM	@�            �@������������������������       ����>9@
           `z@������������������������       ����kӧ	@�           h�@                          �8@.���@            �G@������������������������       ����v/@             @@������������������������       ���n��S@             .@                          �5@ݓ>ț�@�           8�@                            �?��W�q@�           ��@������������������������       �/�7�-@]             c@������������������������       ����!�@7           �@                          �<@L,|��@           �{@������������������������       �a?��\@�            pv@������������������������       ��ax:�7@/            �T@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@      r@     x�@      ?@     �I@     p}@      S@     ��@     �l@     (�@     �v@      :@      �?     @S@      e@      @       @      \@       @     0{@      C@     0r@     �U@              �?     �K@     �R@       @      @      O@      @     �X@      7@      ]@     �G@              �?      1@      <@                      7@              F@      @      N@      (@                      @      2@                      "@              ;@       @     �D@       @              �?      ,@      $@                      ,@              1@      �?      3@      @                      C@      G@       @      @     �C@      @     �K@      4@      L@     �A@                      1@      6@       @      @      9@      @      ?@      &@      4@      2@                      5@      8@              �?      ,@              8@      "@      B@      1@                      6@     �W@      �?      @      I@      @      u@      .@     �e@     �C@                      �?      3@      �?       @      3@      @     �Y@             �A@      (@                      �?      1@      �?       @      ,@              Y@              ?@      (@                               @                      @      @       @              @                              5@      S@               @      ?@             @m@      .@     �a@      ;@                      3@     @R@               @      ?@              m@      &@     `a@      8@                       @      @                                      �?      @      �?      @              5@     �j@     `x@      <@     �E@     pv@      Q@     H�@     �g@     �@     pq@      :@      4@     `c@      m@      4@      @@     `o@     �M@     �g@     `d@     �n@      h@      6@      ,@     �b@     �l@      4@      @@     �n@      M@     `g@      c@      n@     �g@      1@      @      @@     @R@      �?      @      G@      @     �S@     �D@     @V@     �H@              "@     �]@     �c@      3@      ;@      i@     �K@     @[@     �[@     �b@     �a@      1@      @      @      @                      @      �?       @      &@      @      @      @      @       @      �?                      @               @      "@      �?      �?      @              @       @                              �?               @      @       @              �?      M@     �c@       @      &@      [@      "@     �t@      <@     �r@     �U@      @              7@     @Y@      �?      @     �G@      @     �l@      *@     `g@     �F@       @               @      9@               @      @             @Q@      @     �B@       @                      5@      S@      �?      @     �E@      @      d@      @     �b@     �B@       @      �?     �A@      L@      @      @     �N@      @     �Y@      .@     @\@     �D@       @      �?      ;@      G@      @      @     �C@      @      X@      ,@     �V@      >@       @               @      $@      �?       @      6@              @      �?      6@      &@        �t�bub��     hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJƘ�	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Xx��%2@�	           ��@       	                   �;@`vx�V	@�           ��@                            �?�JD��@H           |�@                           �?�cn �@�            Pz@������������������������       ����^��@O            @a@������������������������       ��3��ž@�            �q@                           �?t���@M           Ѝ@������������������������       �3j�Jl@�            pv@������������������������       ����9	@m           ��@
                           �?� qo�	@�            �p@                           �?�U�R@6            @V@������������������������       ���z�W@             F@������������������������       ����!lO@            �F@                           @_�,~%C@p            `f@������������������������       �X����@3             U@������������������������       ��7-�g@=            �W@                          �2@*��k>�@�           ��@                           @���]@�           p�@                          �1@��Neռ@�            0r@������������������������       �*��@x            `f@������������������������       �*��OV@@             \@                           �?���� @           �x@������������������������       ��kH�&��?y             g@������������������������       ������D@�            `j@                           @��@�           ��@                           @}?eG�@
           �y@������������������������       �[�di�#@�             r@������������������������       �h*�F�@H            �_@                           @W#��-�@�           D�@������������������������       �''�40@�           @�@������������������������       �(�}nU@�            �x@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     �s@     �@      4@      K@     �}@      Q@     �@     �k@     ��@     px@      <@      1@     �e@     �k@      .@     �C@     @p@     �E@     �k@     �`@     �p@      m@      2@       @     @a@     �g@      .@      >@     �l@      =@     �i@      Z@     �n@     �d@      ,@             �K@     �N@      �?      &@     �Q@      $@      N@      ?@     �T@     �@@      @              ,@      ?@                      &@             �@@      @     �C@      @                     �D@      >@      �?      &@      N@      $@      ;@      <@      F@      :@      @       @     �T@      `@      ,@      3@      d@      3@     @b@     @R@     �d@     ``@      "@       @      ;@      I@      �?       @     �K@      @     �R@      4@     �P@      I@       @      @      L@     �S@      *@      &@     @Z@      0@     �Q@     �J@     �X@     @T@      @      "@     �A@      ?@              "@      =@      ,@      1@      >@      6@      Q@      @      @      0@      ,@              @      @              @      @       @      4@      �?      @      @      *@              @       @              �?      @       @      $@              @      (@      �?              @      @              @       @      @      $@      �?       @      3@      1@               @      8@      ,@      (@      8@      ,@      H@      @       @      @       @                      $@      @      @      $@      @      >@       @              ,@      "@               @      ,@      $@      @      ,@       @      2@      �?       @     �a@     0r@      @      .@      k@      9@     �@     �U@      �@     �c@      $@              =@     �S@      �?      @     �B@      @     `s@      1@     `d@     �B@      �?              0@      C@               @      2@      @     @^@      &@     �L@      7@                      @      8@                       @             @S@      @     �E@      .@                      &@      ,@               @      $@      @      F@      @      ,@       @                      *@     �D@      �?      @      3@             �g@      @     �Z@      ,@      �?              @      ,@                      $@              \@      �?     �A@      @      �?               @      ;@      �?      @      "@             @S@      @     �Q@       @               @     �[@     �j@      @       @     �f@      4@     �|@     �Q@     x@     �^@      "@              E@      J@               @     �K@      &@      W@      @@     �V@     �B@       @              @@      A@               @      D@       @     �P@      0@     �J@     �A@       @              $@      2@                      .@      @      :@      0@     �B@       @               @     @Q@      d@      @      @     @_@      "@     w@      C@     pr@     @U@      @       @      D@      Z@              @      S@      @      q@      8@      h@      I@      @              =@      L@      @      @     �H@      @     �W@      ,@     �Y@     �A@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���phG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�:H�H:@�	           ��@       	                    �?�I�a�@_           ��@                          �;@>H-C[	@�           �@                          �6@uB���@N           ��@������������������������       ����1�@&           `�@������������������������       ���h.J�@(            {@                           �?�SP��	@�            �p@������������������������       ���z�;�@0            @T@������������������������       ��YL��
@o            �f@
                          �=@D~z���@r           ��@                          �5@<~��I@^           p�@������������������������       �Xu���@�             u@������������������������       �({ӟ5@�            �k@                           �?ʰ)�f@            �A@������������������������       ��ɼdg��?             2@������������������������       �v-�q&x@	             1@                          �3@h<�r�@W           ț@                           @'e/�l@�           P�@                           @	�C�( @�             w@������������������������       ��R�����?F            @Z@������������������������       ����?�4�?�            �p@                           �?7n�!�@�            �y@������������������������       �N@�2�i@             j@������������������������       ��P�k�#@�            �h@                           @�=܆!t@d           @�@                           @��Y��@�           ��@������������������������       �A�(t�\@           @}@������������������������       ��;�
@x            `h@                           �?E�5�v~@�            u@������������������������       �w^!�p�@^            @b@������������������������       ��~0�\�@t            �g@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     �r@     �@      ?@     @P@     0{@     �P@     ��@     �h@     �@      w@      ?@      6@      l@     @s@      2@      I@     Pr@     �G@      v@     �c@     �w@     Pp@      7@      6@     @e@     �l@      1@     �E@     �k@      C@     �i@     �^@     �o@     @h@      6@      "@      b@     @h@      ,@      =@      g@      9@      h@      [@     �k@     @a@      4@       @     @X@     �\@      "@      5@      Z@      3@     `c@      N@     �c@     @W@      @      �?     �G@      T@      @       @      T@      @      C@      H@     �N@     �F@      .@      *@      :@     �B@      @      ,@     �B@      *@      *@      .@     �A@      L@       @      @      @      $@      �?       @      *@              @      @      ,@      4@              $@      4@      ;@       @      (@      8@      *@      @      $@      5@      B@       @              K@     @S@      �?      @      R@      "@     @b@      B@     �^@     �P@      �?              I@      R@      �?      @      N@       @     �a@      =@     �^@     �P@                      2@      G@      �?      @      ?@      @     @Y@      1@     �S@      ?@                      @@      :@                      =@       @     �D@      (@      F@      B@                      @      @              �?      (@      �?      @      @                      �?              �?      �?              �?      @                      @                      �?              @      @                      @      �?      @                                             �S@     �m@      *@      .@     �a@      3@     ��@      C@     �|@     @[@       @              6@     �U@      @       @     �F@      �?     �u@       @     �j@      C@      �?              ,@      >@              @      1@      �?     �h@      @     �V@      (@      �?              @      1@                      �?      �?     �J@              5@      @                      @      *@              @      0@             �a@      @     @Q@      @      �?               @      L@      @      @      <@             @c@      @     @_@      :@                      @      ?@       @      �?      5@              U@      @      I@      ,@                      @      9@       @      @      @             �Q@             �R@      (@                     �L@     �b@      "@      @     @X@      2@     ps@      >@     @n@     �Q@      @              A@     �W@       @       @     �Q@      @     @m@      ,@      e@      A@      @              "@     �Q@               @     �J@      @     �e@      "@     @`@      1@                      9@      8@       @              1@       @      N@      @      C@      1@      @              7@     �L@      @      @      ;@      (@     @S@      0@     �R@     �B@       @              @      4@      @      @      &@      @      E@      @      @@      0@                      1@     �B@      @      �?      0@      @     �A@      &@      E@      5@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�o�>hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?e$h�g@�	           ��@       	                   �5@�tD3�l@�           ,�@                          �2@QV�{�@�           @�@                           �?v=xob@           �y@������������������������       �K��1@R            �_@������������������������       ��Y����?�            �q@                           �?Q1B���@�            �t@������������������������       �L��>,@u            �h@������������������������       ��g��	@\            �`@
                          �<@�(/`+h@%           0~@                          �8@h�C��)@�            Px@������������������������       ��SO�@@�            `l@������������������������       �g�z|�@g            @d@                          @@@[��R`G@9            �W@������������������������       �w�?��@+            @R@������������������������       ���=@             5@                           @��u\~O@�           ��@                          �5@<����	@�           ��@                           �?���IA�@�           (�@������������������������       �p��U��@6           @������������������������       ��D7�::@�            �j@                           �?β�|�	@�           ��@������������������������       ��c>��@�            �h@������������������������       �kM��
�	@s           ��@                          �7@��sw<@�           t�@                           @ol��X"@           ��@������������������������       �"B��j@�           �@������������������������       �z�eW+k@z            @j@                          �:@�0��Q@�            �r@������������������������       �3i�&E	@m            `d@������������������������       �Sy�}�.@\            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        :@      t@     �@      5@     �P@     �|@      T@     �@     @j@     ��@     �v@      B@      �?     �T@     �b@       @      4@      [@      @     �}@      E@     �p@     �Q@      $@             �@@      V@              &@      G@             pu@      8@     �c@      A@      @              1@      C@              @      ?@             �k@      "@     @R@      .@      @              @      4@              �?      2@             �G@      @      3@      "@                      &@      2@              @      *@             �e@       @      K@      @      @              0@      I@              @      .@             @^@      .@     @U@      3@      @              @      6@              @      &@             @T@      (@      E@      *@      @              "@      <@                      @              D@      @     �E@      @              �?     �H@      N@       @      "@      O@      @      `@      2@     �[@      B@      @      �?     �D@     �F@       @       @      J@      @     �\@      $@     �X@      2@       @              ?@      :@       @              9@      �?     �O@       @     @P@      &@      �?      �?      $@      3@               @      ;@       @      J@       @     �@@      @      �?               @      .@              @      $@      �?      ,@       @      (@      2@      �?              @      &@              @      @              ,@      @      &@      0@      �?              @      @              @      @      �?              �?      �?       @              9@     �m@     `v@      3@     �G@      v@      S@     h�@      e@     X�@     pr@      :@      6@     `c@     �j@      *@     �C@      n@      N@      h@     @a@     `k@     �g@      7@      *@      I@     �T@      @      2@     �_@      2@     @^@      K@     @`@      V@      @      *@      E@     �H@      @      .@     �U@      (@     @Q@      >@     @W@     �S@      @               @     �@@              @     �C@      @      J@      8@     �B@      $@              "@     @Z@     �`@      "@      5@     �\@      E@      R@      U@     @V@      Y@      2@              0@      =@      @       @     �@@      @      B@      4@      1@      >@      @      "@     @V@     �Y@      @      *@     �T@     �C@      B@      P@      R@     �Q@      ,@      @     �T@      b@      @       @     @\@      0@     �v@      >@      s@     �Z@      @             �K@     �[@      @      @     @Q@      ,@      s@      *@     �m@     �Q@      �?              C@     �T@       @             �I@      "@     `o@      *@     @f@     �G@      �?              1@      <@       @      @      2@      @     �J@              M@      8@              @      <@     �@@       @      @      F@       @      N@      1@      Q@      B@       @      @      @      .@      �?       @      3@       @     �A@      (@      F@      7@       @              7@      2@      �?      �?      9@              9@      @      8@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJKw�hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @G�1@�	           ��@       	                   �4@���$�@�           J�@                          �2@Z8b(%@K           ��@                           @����O�@?           �@������������������������       ��_����@�            �x@������������������������       ���*1@@             [@                           �?Pw$Z�@           �y@������������������������       ����v@P            �_@������������������������       ��+V�|S@�            �q@
                            �?BeL��5	@B           <�@                           �?GR�i$q	@�            x@������������������������       �R���n@A            @Z@������������������������       �,H[6�	
@�            �q@                           �?���e�@S           p�@������������������������       ��'t	@�            �v@������������������������       ��ۏH�i@j            �@                           �?i�>W�@-           ��@                            �?�>MN܃@j           X�@                            �?n���@�            �t@������������������������       �:_�g���?W            �a@������������������������       ��Aq��@u            @g@                          �0@���s!��?�            0p@������������������������       �
߈�][�?             6@������������������������       �[K�v���?�            �m@                           @A~��J@�           d�@                          �<@u�>���@            X�@������������������������       ��7�_Hi@�            �@������������������������       �m<�~@            �C@                          �5@� 2Ǻ@�            �r@������������������������       �&T���"@k            �e@������������������������       �8/ar@X            @`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �q@     P�@      <@     �J@     �}@      U@     Џ@      l@     H�@     �w@      5@      *@     @i@     �u@      4@     �E@     �t@     �N@     px@      g@     �u@      p@      0@      @     �O@     �_@       @      (@     ``@      *@     @n@     �P@     `c@     �X@       @      @      >@     �Q@              @      M@      @     �c@     �B@     �U@     �I@      �?              3@      I@              �?      H@      �?     ``@      <@     �R@      F@              @      &@      5@              @      $@       @      ;@      "@      *@      @      �?       @     �@@     �K@       @       @     @R@      $@      U@      >@      Q@      H@      �?              0@      .@                      1@      �?      B@      "@      9@       @               @      1@      D@       @       @      L@      "@      H@      5@     �E@      D@      �?      @     `a@     �k@      2@      ?@      i@      H@     �b@     @]@     �g@     �c@      ,@      @      ?@     �P@      @      ,@     @Q@      2@     �G@     �C@     �K@     �@@      @      �?      "@      2@                      8@      @      1@      @      :@       @              @      6@      H@      @      ,@     �F@      .@      >@      A@      =@      ?@      @      @      [@     `c@      .@      1@     �`@      >@     �Y@     �S@      a@     �_@       @      �?      G@     �N@      $@      $@     �E@      3@      A@      :@      J@     �L@      @       @      O@     �W@      @      @     @V@      &@      Q@      J@      U@     @Q@      @      �?      U@     �i@       @      $@     �a@      7@     ��@      D@     �z@     @^@      @              3@     �P@       @      @      ;@       @     �q@      *@     �a@      9@                       @     �E@       @      �?      4@       @     �a@      @      T@      5@                              3@       @              @      @     �S@              8@       @                       @      8@              �?      *@      @     �O@      @      L@      *@                      &@      7@               @      @             �a@      "@      O@      @                              �?                      @              1@                      �?                      &@      6@               @      @              _@      "@      O@      @              �?     @P@     �a@      @      @      ]@      .@     �u@      ;@     r@      X@      @      �?      E@      Y@       @      @     @S@      @     �r@      &@     `h@      Q@      @      �?      B@     �W@       @      �?     �P@      @     �r@      &@     �g@     @P@      @              @      @               @      &@              @              @      @                      7@     �D@      @      @     �C@      "@      E@      0@     �W@      <@       @              @      ;@      �?      �?      8@      �?      A@      @     �O@      &@       @              2@      ,@      @      @      .@       @       @      *@      ?@      1@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJrg�5hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?[�v?=9@�	           ��@       	                    �?��ҿu@           ��@                           �?����@(           @}@                          �<@!�wB<@h            `e@������������������������       ��y�z|{@]            �b@������������������������       ��k�d�?             5@                           �? ͬ%j@�            �r@������������������������       ��+z���@^            `b@������������������������       �����U@b            �b@
                          �=@'���q�@�           ��@                          �1@fr/dz@�           ��@������������������������       ���u�P�?~            �i@������������������������       ���B��@Z           @�@                            �?XЈq	@             >@������������������������       ��(;��e@             3@������������������������       �=*,I�R @             &@                           @w��c,@}           Ƥ@                           �?�6_��	@�           ��@                           �?:����	@�           t�@������������������������       �3|[�%t	@�            �y@������������������������       ��g���	@�           �@                            �?��I�@�            y@������������������������       �����@F            �Z@������������������������       ���t|�@�            `r@                          �8@��^��@�           ԑ@                           @�M؟�@4            �@������������������������       �{p��3�@+           ��@������������������������       ��E�g@	             &@                           @��5ܘ@�            �n@������������������������       ��y�~�@�            @m@������������������������       ��7���� @             &@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �s@     ��@      @@     �F@     `x@     �U@     ��@     �l@     p�@     0v@      9@       @      X@     �f@      �?      @     �W@      ,@     }@      D@     �p@     @U@      @       @     �L@      U@      �?      @     �L@      @     �Y@      :@     @T@     �G@      �?       @      ,@      >@                      5@              L@       @      :@      ,@               @      (@      3@                      3@              L@       @      9@      "@                       @      &@                       @                              �?      @                     �E@      K@      �?      @      B@      @     �G@      2@     �K@     �@@      �?              7@      8@      �?      @      1@      @      :@      (@      2@      0@      �?              4@      >@                      3@              5@      @     �B@      1@                     �C@     @X@                     �B@      $@     �v@      ,@      g@      C@      @              C@     @X@                     �@@      "@     �u@      &@     �f@     �A@      �?              @      1@                      ,@             �^@      �?     �A@      @      �?              @@      T@                      3@      "@     �l@      $@     @b@      <@                      �?                              @      �?      &@      @      @      @      @                                               @      �?      @      @       @      �?      @              �?                               @              @              �?       @              7@     �k@     �w@      ?@      D@     �r@      R@     ��@     �g@     (�@     �p@      3@      7@     �b@      l@      8@      >@      j@      K@     �k@     �d@      k@     �f@      1@      7@     @]@     @c@      6@      5@     �b@     �F@     ``@     �_@     �d@     �b@      0@      ,@      >@     @R@      .@       @     �O@      (@      H@      K@     �D@      L@      @      "@     �U@     @T@      @      3@     @U@     �@@     �T@      R@     �^@     �W@      *@              ?@     �Q@       @      "@      N@      "@      W@     �D@     �J@      @@      �?              &@      .@              @      *@      @     �C@      @      (@      @      �?              4@      L@       @      @     �G@      @     �J@      C@     �D@      9@                     �R@     �c@      @      $@      V@      2@     `w@      8@     �r@      V@       @             �J@     @]@      @      @     �N@      .@     �t@      0@     �m@     �L@       @              J@      ]@      @       @     �L@      *@     �t@      0@     �m@      L@       @              �?      �?              �?      @       @                      �?      �?                      5@     �C@      �?      @      ;@      @     �F@       @     �O@      ?@                      1@     �B@      �?      @      :@             �F@       @      O@      ?@                      @       @                      �?      @                      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ$�YhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �4@���%:Y@�	           ��@       	                    �?kl%ڱ@�           \�@                           �?��:�.@�           0�@                           �?j���g@�            �h@������������������������       ��Ǵ���@1             S@������������������������       ��kd��@Q             ^@                           �?��t���?4            ~@������������������������       �-�. @�             p@������������������������       ������o�?�             l@
                           @�`�v\W@�           đ@                           @{n1���@l           ��@������������������������       ��̠z�\@�            x@������������������������       �M G��@w            �g@                          �3@�&��[@k           ��@������������������������       ����\�@#           �{@������������������������       ��ۄ��9@H            @^@                           @
3�@Z�@8           d�@                           �?�"j�*l	@C           t�@                           �?ES1<#�@�            �u@������������������������       ��Jbp�@�            Pp@������������������������       �c���C@:             U@                          �:@�__]�	@g            �@������������������������       ��^��Z	@�           ��@������������������������       ���	��	@�            �r@                           �?)��8@�           ��@                           @w���!�@�            �v@������������������������       ��vҿ@�            Pq@������������������������       �����_�@8            @V@                           @�%D�.@           pz@������������������������       �-�y	@�            Pw@������������������������       �Cv�D	@!             I@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@     Pr@     ��@      @@     �N@      @     �P@     ��@      m@     Ї@     Pu@      @@      @     �X@     �n@      @      3@     �f@      (@     Ѓ@     �W@     �w@     �`@      @              >@     �R@              @     �H@      @      t@      ;@     �a@      8@                      &@     �B@              �?      9@      @      I@      2@     �B@      (@                       @      *@                      $@              6@      �?      6@      @                      "@      8@              �?      .@      @      <@      1@      .@      @                      3@      C@              @      8@              q@      "@     �Y@      (@                      "@      5@              @      3@             @b@      @     �F@      @                      $@      1@                      @             �_@       @      M@      @              @      Q@     �e@      @      *@     �`@      @     �s@     �P@     �m@     �[@      @      @     �B@      W@      @       @     �X@      @     @Z@     �L@     @V@     �Q@      @      @      9@     �O@      @      @     @S@      @     �N@      ;@     �P@     �I@              �?      (@      =@              @      6@      �?      F@      >@      7@      4@      @              ?@      T@       @      @      A@      @     �i@      $@     �b@      D@                      3@     �P@       @      @      =@             @d@      @     �_@      9@                      (@      *@                      @      @     �F@      @      8@      .@              ,@     `h@     �s@      :@      E@     �s@     �K@     �w@     @a@     �w@     �i@      <@      ,@     `b@     @j@      5@      B@     @k@     �@@      e@     �Z@     �f@     �b@      5@             �G@      K@      @      @     �I@      �?     �Q@      4@      H@     �B@      @              E@      F@      @      @     �F@      �?      B@      *@      B@      >@      @              @      $@                      @             �A@      @      (@      @       @      ,@      Y@     �c@      2@      >@     �d@      @@     �X@     �U@     �`@     @\@      ,@      @     �R@      ]@      "@      :@     �[@      3@     @R@      M@     �Y@     �M@      $@      "@      9@      D@      "@      @      L@      *@      9@      =@      @@      K@      @              H@     �Z@      @      @     �X@      6@     @j@      ?@      i@      L@      @              =@      N@              @     �M@      &@     �X@      "@     �S@      0@       @              4@     �G@               @      A@      @     �U@      @     �O@      &@                      "@      *@              �?      9@      @      (@       @      0@      @       @              3@      G@      @      @     �C@      &@      \@      6@     @^@      D@      @              &@      E@      @      @     �@@      "@     �Z@      4@     @\@     �@@                       @      @       @              @       @      @       @       @      @      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ �u)hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @b��.�2@�	           ��@       	                    �?�zˋ7�@?           ��@                           �?��qp �@�           P�@                          �8@�d|��'@�            �s@������������������������       �mfA�W@�            �m@������������������������       �p����G@0            @T@                            �?:��ln@�            �t@������������������������       ��.$i�@             i@������������������������       ����*CF@Q            @`@
                          �3@V�O�~|	@�           $�@                           �?AI�u��@           `z@������������������������       �%�1��@�            Pq@������������������������       ���K�6@^             b@                            �?n�QW�	@�           ��@������������������������       �: ?TɈ	@�            �r@������������������������       ��/P�Y�	@�           ��@                           @��?a�@a           ؛@                           �?���U�@	           ��@                           �?.���@           �}@������������������������       ������5@�             q@������������������������       ��,f{ @}             i@                           @�ڐ��-@�           x�@������������������������       �����@�           ��@������������������������       �:Qꎳ�@             3@                          �6@� ~��@X           x�@                           �?X����@�            @t@������������������������       ������@q            �d@������������������������       �΀{�`�@f            �c@                           @��5�	@�            `i@������������������������       ���ϔ��@_            @b@������������������������       ����X@"            �L@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     �q@     �@      5@     �J@     �}@     @T@     (�@     `j@     ��@     �w@      8@      8@      i@     �s@      1@     �D@     `s@      O@     �u@     �f@     Pv@     p@      5@      �?      N@      T@       @      @      U@      @     @b@      >@      d@     �Q@      @      �?      >@      A@       @      @     �A@      @     �T@      4@     �N@     �D@                      6@      9@       @      @      9@      @     �R@      (@      G@      6@              �?       @      "@              @      $@               @       @      .@      3@                      >@      G@                     �H@             �O@      $@     �X@      >@      @              ,@      :@                      7@              @@      @     �S@      4@      @              0@      4@                      :@              ?@      @      5@      $@              7@     �a@     �m@      .@      A@     @l@     �L@      i@     �b@     �h@     @g@      1@      @      A@      O@              @     �I@      @     @W@     �H@     �O@     �H@      @      @      ?@      A@              @     �B@      @      I@      @@      C@     �B@      @              @      <@               @      ,@      �?     �E@      1@      9@      (@              2@     �Z@     �e@      .@      <@     �e@     �I@     �Z@     @Y@     �`@      a@      *@      �?     �@@      F@      @      ,@      E@      *@      G@      7@     �A@     �D@      @      1@     @R@     @`@      &@      ,@     �`@      C@     �N@     �S@     �X@      X@      $@      �?     �T@     �l@      @      (@     �d@      3@     X�@      ?@     �|@     �^@      @      �?      L@     �b@      @      �?     �X@      *@     `�@      3@      t@      Q@       @      �?      7@      M@                      7@       @      l@      @     @]@      $@              �?      ,@     �A@                      1@      �?     @_@      @      Q@      @                      "@      7@                      @      @      Y@      @     �H@      @                     �@@     �V@      @      �?      S@      @     �r@      (@     `i@      M@       @              @@     �V@       @      �?     @R@       @     �r@      $@     �h@     �K@       @              �?              �?              @      @       @       @      @      @                      ;@      T@      �?      &@     @P@      @     �_@      (@     �a@     �K@      �?              2@      H@      �?      @      A@      �?     �Y@      @      T@      <@      �?               @      8@      �?      @      5@      �?      K@       @      A@      1@                      $@      8@              �?      *@             �H@       @      G@      &@      �?              "@      @@              @      ?@      @      8@       @      O@      ;@                      @      <@              @      ,@      @      0@      @     �H@      3@                      @      @                      1@               @      �?      *@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��3hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�<@`�U@�	           ��@       	                     �?oY:�_f	@�           ��@                           �?���i	@9           �}@                           �?\u=t@x             g@������������������������       �(�nb��@+            @Q@������������������������       �[h�2G@M            �\@                           �?�ɥF]	@�            0r@������������������������       ����@7            @W@������������������������       ��ӟ��	@�            �h@
                           �?�:W	@�           0�@                           @O���@	           �y@������������������������       �Y��@x            �g@������������������������       ��^ۨ�!@�            �k@                            �?�!#�>�	@�           ��@������������������������       ��!Z��H
@u            �f@������������������������       ������E	@?           �@                           �?[nF��@�           D�@                            �?QR��X�@�           0�@                           �?�b`@/��?s             g@������������������������       ��u�M�?=            @W@������������������������       ��n�*G�?6            �V@                           @�t�:�@u           p�@������������������������       �u�o^�@�            �v@������������������������       �
��׻I@�             l@                          �4@��/�@�           p�@                           @ ��S@�           ؈@������������������������       �U��4\f@�           ��@������������������������       ��[��]�@T            �`@                            @|��3_d@�           �@������������������������       �����e@}           P�@������������������������       �8����@b            �b@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        ,@     �r@     P�@      6@     �K@     �|@     �W@      �@      k@     ��@     �v@     �A@      (@     �d@     @k@      1@     �A@     @o@      N@     �j@     @`@     0p@      g@      @@      @     �I@     �P@      @      "@     �Q@      4@     �M@      F@     �U@     �G@      ,@      @      *@      9@              @      ?@      @     �@@      ,@      C@      (@       @      @       @      $@                      ,@      @      (@      &@      $@       @      �?              &@      .@              @      1@       @      5@      @      <@      $@      �?      �?      C@      E@      @       @     �C@      ,@      :@      >@     �H@     �A@      (@              $@      0@                      *@      �?      2@      @      7@      "@              �?      <@      :@      @       @      :@      *@       @      ;@      :@      :@      (@       @     �\@     �b@      ,@      :@     �f@      D@      c@     �U@     �e@     @a@      2@              ;@     �M@       @      @     @P@      "@     �T@      >@     @S@      G@      @              *@      8@       @              4@       @     �H@      .@     �F@       @      @              ,@     �A@              @     �F@      �?      A@      .@      @@      C@       @       @     �U@      W@      (@      4@     �\@      ?@     �Q@      L@     �W@      W@      (@       @      9@      0@      @      (@      3@      "@      .@      6@      4@      @@      �?      @      O@      S@      @       @      X@      6@     �K@      A@     �R@      N@      &@       @     @a@      u@      @      4@     `j@     �A@     ��@     �U@     ��@      f@      @             �@@      Z@               @     �E@      @     �u@      5@     @f@     �C@                      �?      $@                      "@      �?      Z@      @      H@      @                              @                      @              N@              3@       @                      �?      @                       @      �?      F@      @      =@      @                      @@     �W@               @      A@      @     �n@      0@     @`@     �@@                      :@     �G@                      2@      @     �e@      "@     �R@      0@                      @     �G@               @      0@             @R@      @      L@      1@               @     @Z@      m@      @      2@      e@      >@     0{@     �P@     �v@     @a@      @             �C@     �^@      @      @     �P@      @     0r@      =@     �f@     �J@                      ;@     �Y@              @     �H@      @     �o@      =@     �b@     �E@                      (@      3@      @      @      1@      @     �B@              =@      $@               @     �P@     �[@       @      (@     �Y@      8@      b@     �B@     �f@     @U@      @       @      K@     �W@      �?      (@     �U@      7@     @Z@      <@     @c@      L@       @              (@      .@      �?              0@      �?     �C@      "@      <@      =@      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJu�+hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?Ôvg"\@�	           ��@       	                   �2@Ҋ��^w	@�           d�@                            @mfo��N@�            �t@                           �?oŢ��Q@i             f@������������������������       ���89@6            @V@������������������������       �c�1�R�@3             V@                           @k@�R@]            @c@������������������������       �2��}o�@2            �T@������������������������       �Z�_�[@+             R@
                           �?Z��	@0           8�@                           �?:@D��@�            �u@������������������������       �}A�uW�@T            @^@������������������������       �A���14@�            `l@                           �?��؉�Y
@M           ��@������������������������       ����K[N	@�            �r@������������������������       ��l��[
@�            �@                          �7@(61Թ�@�           �@                           �?yO�@Z            �@                          �1@x#	�� @~            �@������������������������       �m� (:�?t            `g@������������������������       ��^�?@
           �z@                           @-9�$��@�           ��@������������������������       �u��^�7@4           �~@������������������������       ��,J_o�@�           ȃ@                           @X,���@`           @�@                           �?F0���@c            �c@������������������������       ��4���@/            �Q@������������������������       ��{�j$@4             V@                          �<@_-���<@�            �x@������������������������       ��{�1�@�            �s@������������������������       ���&� �@1            @S@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     v@      �@      B@     �F@     �{@     �U@     X�@     �g@     ��@     @v@     �A@      3@     �i@     �p@      :@     �@@     �j@      J@     �l@      _@     �n@     �f@      =@       @      C@      I@      �?      @      E@             �S@      :@      K@      =@      @              1@      4@                      ;@              G@      1@      <@      3@      @              @      @                      &@              >@      (@      .@      *@                      (@      1@                      0@              0@      @      *@      @      @       @      5@      >@      �?      @      .@             �@@      "@      :@      $@               @      "@      0@              �?      @              :@      @      *@      @                      (@      ,@      �?      @      &@              @      @      *@      @              1@     �d@     �k@      9@      :@     �e@      J@     �b@     �X@     �g@     �b@      :@              G@     @Q@       @      @      H@      �?     �M@      (@     @R@      ?@       @              0@      4@                      *@              >@       @      =@      &@                      >@     �H@       @      @     �A@      �?      =@      $@      F@      4@       @      1@     @^@      c@      7@      5@      _@     �I@     �V@     �U@     @]@      ^@      8@      @      5@      K@      @      &@      L@      (@     �F@      2@     �D@      ?@      @      ,@      Y@     �X@      2@      $@      Q@     �C@     �F@      Q@      S@     @V@      3@      �?     �b@     Ps@      $@      (@     @l@     �A@     ��@     �P@     ~@      f@      @             @X@     `o@      $@      @     �b@      6@     ��@      9@     �v@     @]@      @             �@@     @P@              �?      F@             �r@       @     `a@      7@       @              @      &@              �?      &@              [@      �?     �G@      @       @              >@      K@                     �@@             `h@      �?      W@      4@                      P@     @g@      $@      @     �Z@      6@     Px@      7@     �k@     �W@       @             �@@     @W@      @      @     �G@      2@     �c@      2@     �P@      I@       @              ?@     @W@      @      @      N@      @      m@      @     @c@      F@              �?     �I@      M@              @     �R@      *@     �_@     �D@     @^@     �M@       @              3@      4@                      0@      @      =@      4@      6@      8@      �?               @      @                      @              ,@      "@      $@      1@                      &@      .@                      "@      @      .@      &@      (@      @      �?      �?      @@      C@              @     �M@      @     @X@      5@     �X@     �A@      �?      �?      1@      ?@              @      D@      @     �U@      2@     �V@      6@      �?              .@      @                      3@      �?      $@      @      "@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ'�f	hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@���1e@�	           ��@       	                    �?�
ɓf�@k           �@                            �?2<���P@�           ��@                           �?Ib"X�� @�             k@������������������������       ��a�s���?B            �Z@������������������������       ��`���! @G            �[@                           @z����@f           0�@������������������������       �o)�7@�            `q@������������������������       ��`w �O @�             s@
                           @�	9��@|           ��@                           �?���a�O@J           8�@������������������������       �-�C�<@�            �s@������������������������       �BL�M �@t           X�@                           �?[� 9�@2           p~@������������������������       ��(L���@z            �g@������������������������       ���rM�@�            �r@                           @���-�@7           �@                           �?wg��~	@�           �@                          �<@D���l@�            �p@������������������������       ���dYR@�            �h@������������������������       ���G3@+            �P@                           �?�����	@           ��@������������������������       ��8�n�	@�            �r@������������������������       �b�e���	@J           ��@                           @�Dz��v@�           ��@                          �7@e51�p@�            @y@������������������������       �Zz�1j@i            �c@������������������������       ��V�2%@�            �n@                           �?�}|@�             l@������������������������       �)�Ύ�(@3            �U@������������������������       ��0w4[1@U            `a@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     `r@     �@      @@     �M@     �{@     �V@     `�@     �k@     ��@     �x@      7@      @      _@     0r@      @      A@     @k@      B@     ��@     �Y@     �~@     @e@      &@              F@      [@      �?      "@     �M@       @     �t@      5@     �e@      G@      @              @     �@@              �?      @             �V@       @      P@      (@                               @              �?      @             �I@       @      @@      @                      @      9@                                      D@              @@      @                     �B@     �R@      �?       @      J@       @     @n@      3@     @[@      A@      @              =@      :@      �?      @      @@       @     �V@      0@      F@      ?@       @               @     �H@              @      4@             �b@      @     @P@      @      �?      @      T@     �f@      @      9@     �c@      A@      w@     @T@     �s@      _@       @      @      J@     @]@      @      ,@      Z@      1@     �m@     �C@     @l@      V@      �?      @      >@     �C@      �?      @     �G@      @     �G@      7@     @P@     �G@      �?              6@     �S@      @       @     �L@      $@     �g@      0@      d@     �D@               @      <@     �P@      �?      &@     �K@      1@     �`@      E@     @V@      B@      @       @      $@      ?@              $@      *@      "@     �J@      4@      6@      1@      �?              2@     �A@      �?      �?      E@       @      T@      6@     �P@      3@      @      *@     @e@     �o@      9@      9@     `l@     �K@     �r@      ^@     �r@     @l@      (@      *@     �^@     �f@      1@      6@      d@     �H@     @]@     @X@     @a@     �d@      (@              ?@      @@               @      H@      @      E@      2@     �G@      D@      �?              9@      <@                     �@@      @     �C@       @     �D@      4@      �?              @      @               @      .@              @      $@      @      4@              *@      W@     �b@      1@      4@      \@      G@     �R@     �S@     �V@     @_@      &@      @      <@     �L@      $@       @     �C@      :@      5@      8@     �@@      J@      @      "@      P@     @W@      @      2@     @R@      4@      K@     �K@      M@     @R@      @             �G@      R@       @      @     �P@      @      g@      7@     �c@     �N@                      ?@     �H@                      A@      �?     `b@      "@     �X@     �A@                      $@      7@                      @      �?     �R@       @     �@@      $@                      5@      :@                      =@             @R@      @     @P@      9@                      0@      7@       @      @     �@@      @     �B@      ,@      N@      :@                              @      @              1@              4@      @      9@       @                      0@      1@      @      @      0@      @      1@      @     �A@      2@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ+��_hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�F��@�	           ��@       	                    @L#3B�	@V           �@                          �1@�0�vs[@�           А@                           �?;��0�@�            �q@������������������������       ���@�B@w            �f@������������������������       ��ŕr*�@A             Y@                           �?�����@           ؈@������������������������       ���l��|@�            �o@������������������������       ����ys}@b           ��@
                          �2@�cm9��@�           �@                           @��9�	 @_           `�@������������������������       �x�aa���?�            u@������������������������       ��zŗ{@�            `o@                           �?���c'�@:           P@������������������������       �S��qˉ�?h            `d@������������������������       ���t�$U@�             u@                           @�?.��@Q           P�@                           �?/ϫ�;�	@�           H�@                          �>@I�
p@�            �r@������������������������       �+�x
�i@�            p@������������������������       �<��@            �C@                          �9@k�8&��	@           P�@������������������������       ���{$R	@           P{@������������������������       ���L���	@�            Pw@                           @ڜ��@�           �@                           @r	�N�W@           �|@������������������������       �i���$�@�            �q@������������������������       �Z~r�F�@m            �f@                           @t��6 �@o            `f@������������������������       ��O�ek�@G            @]@������������������������       �,�)Tr�@(             O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@      r@     ��@      :@     �K@      |@     �Q@     8�@     �k@     0�@     v@      ;@      @      \@     �r@      @      <@     @l@      7@     �@      U@     P@     `a@      @      @      S@     `c@      @      7@     �c@      3@     `o@      P@     @l@     @V@      @       @      2@      C@                      =@              X@      2@      L@      8@               @      &@      8@                      :@              J@      $@      C@      2@                      @      ,@                      @              F@       @      2@      @              @      M@     @]@      @      7@     �_@      3@     `c@      G@     @e@     @P@      @              7@     �E@              @      7@      @      O@      (@     @Q@      &@              @     �A@     �R@      @      4@      Z@      *@     @W@      A@     @Y@      K@      @              B@     �a@      �?      @     �Q@      @     `~@      4@     0q@      I@                      1@     @R@      �?      @      :@      �?     �s@      @     @_@      6@                      @      D@                      @      �?     �i@      @     @P@      "@                      *@     �@@      �?      @      3@             �Z@       @      N@      *@                      3@     @Q@              �?      F@      @     �e@      ,@     �b@      <@                      �?      9@                      @             �T@       @      G@       @                      2@      F@              �?     �C@      @     �V@      (@      Z@      :@              &@     @f@     �p@      4@      ;@     �k@     �G@     �r@      a@     s@     �j@      4@      $@     �`@      f@      1@      8@     `b@      B@      `@     @\@      d@     �a@      4@              A@      J@      @      @      C@      �?      M@      (@     �I@     �B@      @              ;@     �H@      @      �?      ?@      �?      L@      @     �G@      A@      @              @      @              @      @               @      @      @      @              $@      Y@      _@      ,@      1@     @[@     �A@     �Q@     @Y@     @[@      Z@      1@       @      L@     @R@      @      ,@     �R@      .@     �B@     �H@      O@     �D@      @       @      F@     �I@       @      @      A@      4@     �@@      J@     �G@     �O@      $@      �?      F@     �V@      @      @     �R@      &@     �e@      7@      b@     @R@              �?      2@     �R@      �?      @      F@      &@      a@      0@     �Z@     �I@              �?      @     �F@               @      5@      @      Y@      @      P@      =@                      *@      =@      �?      �?      7@      @     �B@      "@     �E@      6@                      :@      1@       @              ?@              B@      @      C@      6@                      5@      ,@      �?              5@              @@      �?      2@      "@                      @      @      �?              $@              @      @      4@      *@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�R8hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?@Ü�V@�	           ��@       	                    �?��aZ>	@           @�@                          �;@>�=d��@0           �~@                          �5@Ң���@           P{@������������������������       ����,U@�            Pq@������������������������       �c����@i             d@                          �<@�I4Vu@(             L@������������������������       ��g�L@	             *@������������������������       �,�)g�@            �E@
                          �3@Yv맞�	@�           ��@                           @1���W/@�             r@������������������������       ����Y�@�            `q@������������������������       ��[���@             (@                           �?l�02�
@           �@������������������������       �E�u�]@�             q@������������������������       �����;
@f           x�@                           �?{K�H@�           �@                           @�*��@�           8�@                            �?��`��� @]           h�@������������������������       �A2Ē��@�            �s@������������������������       ��Q���?�            �n@                           �?�BS;
�@�            @k@������������������������       �/�B�op@M            �_@������������������������       �Ύ6My@:             W@                          �4@I�3ɖ0@�           ȗ@                            �?��HԄ�@�           0�@������������������������       �pz�D�@}            �g@������������������������       �NK�h�@u           8�@                           @�3?�@�           `�@������������������������       �����}@�           0�@������������������������       ���9�f@             C@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        1@     �r@     ؁@      5@      L@     �y@     @W@     �@     @m@     ؇@     �w@     �@@      0@     @f@     �n@      (@      =@     �j@     �K@     �n@     `b@      m@     �j@      <@       @      J@     �T@              @      F@      @     �\@      @@      Y@     �K@      �?             �F@     @S@              @     �C@      �?     @[@      ;@     �W@      D@      �?              5@     �B@              @      4@      �?     �U@      1@     �N@      =@      �?              8@      D@              �?      3@              6@      $@     �@@      &@               @      @      @               @      @       @      @      @      @      .@               @      @                              �?       @       @              @                              @      @               @      @              @      @      @      .@              ,@     �_@     �d@      (@      7@     `e@      J@     @`@     �\@     �`@     �c@      ;@      @      ?@     �A@       @              ?@      @     �K@      =@     �E@      I@      @      �?      ?@      A@       @              =@      @     �K@      =@      E@      H@      �?      @              �?                       @      �?                      �?       @       @      $@     �W@      `@      $@      7@     �a@     �F@     �R@     �U@     @V@     �Z@      8@              0@      J@       @      &@      I@      @      C@      4@      B@     �C@      @      $@     �S@     @S@       @      (@     �V@     �D@     �B@     �P@     �J@      Q@      2@      �?     �^@     @t@      "@      ;@      i@      C@     ��@     �U@     ��@     �d@      @              <@     �Y@              @      E@      (@     @w@      ,@     �d@     �@@      @              4@     @Q@                      :@      "@     �q@      @     �]@      5@       @              $@      G@                      3@      @      c@      @      L@      1@       @              $@      7@                      @      @     �`@      �?      O@      @                       @      A@              @      0@      @     �U@       @     �G@      (@      �?              @      6@              @      $@      @      M@      @      *@       @                       @      (@                      @              <@      @      A@      @      �?      �?     �W@     �k@      "@      8@     �c@      :@     �y@     @R@     �v@     �`@       @              :@     @\@      @      @     �J@      "@      r@      <@      h@      L@                      @      9@              �?      ,@      �?     �V@      (@      ;@      ,@                      3@      V@      @      @     �C@       @     �h@      0@     �d@      E@              �?      Q@      [@      @      3@     @Z@      1@     �_@     �F@     �e@     �S@       @      �?      N@      Z@      @      3@     �X@      *@     �^@     �B@     `e@      S@       @               @      @      �?              @      @      @       @       @       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�=;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @-S�]@�	           ��@       	                   �9@�[�r�@g            �@                           �?E؝�H@*           `�@                           �?���7��@�           �@������������������������       �N���0@            |@������������������������       �:b�u	@�           �@                          �2@w`��@D           ��@������������������������       ��qUA@g             e@������������������������       �{Fz �@�            �v@
                           �?�O��
@=           �~@                           @ѕ��r	@y            �g@������������������������       �5�2Ft�@q            �e@������������������������       ���	M�1@             0@                          �;@�
@�            �r@������������������������       �t5��Sp@K            @]@������������������������       �QM>�B{
@y            �f@                          �4@�|�@ @*           $�@                           �?�ڤC{�@A           �@                           @��
D���?�            @x@������������������������       �{��D�?�            �r@������������������������       �˽���}@=            @V@                          �1@x{���<@Y           ��@������������������������       ��>A��@u            �g@������������������������       ����d �@�            0v@                           �?X���@�           0�@                           @b��,�@�            �o@������������������������       �h�9ʙ@E             _@������������������������       �hc^�<@T            @`@                          �8@E�'߱@P           @�@������������������������       ���X���@�            �s@������������������������       �|�j�?�@�            �m@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     �@      @@     �M@      |@      V@     ��@     @j@     ��@     �v@     �@@      .@     @h@      u@      7@     �E@     �s@     @Q@     Pu@     �d@     @x@     �o@      >@       @     `b@     @p@      2@      <@      p@      D@     �r@     @[@     0t@      f@      2@       @     �\@     �g@      .@      9@     `f@      ?@     �d@     @S@      k@     �]@      0@              =@     �T@       @      $@     @R@      "@     @V@      6@     @U@      F@       @       @     �U@     @Z@      *@      .@     �Z@      6@     �S@     �K@     ``@     �R@      ,@              @@      R@      @      @     �S@      "@      a@      @@     �Z@      M@       @              @      9@                      5@              P@      @      B@      (@                      <@     �G@      @      @      M@      "@      R@      9@     �Q@      G@       @      @     �G@     �S@      @      .@     �N@      =@      C@     �K@     @P@      S@      (@      �?      0@      >@       @      @      8@      3@      &@      ,@      5@     �E@       @      �?      .@      >@       @      @      4@      ,@      &@      ,@      3@     �D@                      �?                              @      @                       @       @       @      @      ?@      H@      @       @     �B@      $@      ;@     �D@      F@     �@@      $@              $@      4@                      3@      @      .@      5@      3@      @       @      @      5@      <@      @       @      2@      @      (@      4@      9@      <@       @      �?     �V@     `m@      "@      0@     ``@      3@     ��@      G@     0{@     @\@      @             �A@     �^@      @      @      I@       @     �z@      1@     �k@      D@       @              (@      G@               @      (@              k@      @      V@      @       @              "@      >@                      @             `f@             @Q@      @                      @      0@               @      @             �B@      @      3@               @              7@     @S@      @      @      C@       @     �j@      ,@     �`@     �@@                      @      <@              @      *@              T@      @      I@      @                      4@     �H@      @              9@       @     �`@      &@      U@      :@              �?      L@      \@      @      $@     @T@      1@      j@      =@     �j@     @R@      �?      �?      *@     �K@              �?      (@      (@     �P@      (@     @Q@      (@              �?      &@      >@              �?       @      (@      8@      �?      ?@      @                       @      9@                      @             �E@      &@      C@      @                     �E@     �L@      @      "@     @Q@      @     �a@      1@      b@     �N@      �?              2@      B@       @      @      D@      @     �W@       @      U@      ;@      �?              9@      5@      @      @      =@              G@      .@      N@      A@        �t�bub���      hhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�C�dhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�0�̓a@�	           ��@       	                    �?X{.1	@�           8�@                           �?:7�+@,           �~@                          �:@�%�W��@}            @j@������������������������       �g��_�@i            �e@������������������������       ��n=|i�@             C@                          �4@=����@�            �q@������������������������       �aZ����@K            �_@������������������������       ��0�Js@d            �c@
                          �8@�P0D�	@�           |�@                            @���!�@�           ��@������������������������       ���e�H	@           �y@������������������������       ������@�            �u@                           �?�R?�x
@�            �v@������������������������       ��`��q;@             9@������������������������       �3�&u�M
@�             u@                            @E\8�+/@�           ��@                          �5@Q�N�!@�           ��@                          �4@�fl1�8@�           @�@������������������������       ��ol���@s           ��@������������������������       �t�}V�E@p            `g@                           �?b	�KE@�           p�@������������������������       �8V��.(@v            �f@������������������������       �\}���@=           �@                          �3@}�	I98@           �{@                           @��;��@v             h@������������������������       ��1 E@%             M@������������������������       �U�����?Q            �`@                           @M��(��@�            �o@������������������������       �!��/��@w            �g@������������������������       �6��)�	@)            �O@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        3@      q@     Ѐ@      9@      M@      }@     �T@     (�@     �n@     ��@     �w@      ?@      3@     �c@     �l@      $@     �B@      m@      F@     �l@     �d@     �p@     �h@      9@       @     �G@     �V@              $@     �J@       @     �Z@      >@     @W@      M@      @       @      4@      ;@                      5@              P@      @     �H@      5@      �?              (@      5@                      0@             �L@      @      G@      ,@      �?       @       @      @                      @              @              @      @                      ;@     �O@              $@      @@       @      E@      9@      F@     �B@      @              @      4@                      *@      �?     �@@      $@      7@      5@      �?              7@     �E@              $@      3@      �?      "@      .@      5@      0@       @      1@     �[@     �a@      $@      ;@     `f@      E@      _@      a@     �e@     �a@      5@      $@      T@     �X@      @      0@     `a@      4@     �W@     �R@      ^@     @W@       @      @      H@     �J@      @       @      O@      ,@      O@     �I@     �J@      I@      @      @      @@     �F@      �?       @     @S@      @     �@@      8@     �P@     �E@       @      @      ?@      E@      @      &@      D@      6@      =@     �N@      J@     �G@      *@       @              @                      �?      �?              @              @      @      @      ?@      C@      @      &@     �C@      5@      =@      K@      J@      E@       @             �\@     @s@      .@      5@      m@     �C@     ��@     @T@     ��@      g@      @             @W@     �o@      $@      (@     �h@     �A@     0�@     �N@     �z@     �b@      @             �B@     @e@      @      @     �W@      ,@      |@      5@     �r@      Q@      @             �@@     �`@      @      @     @S@      @     �x@      4@     �n@     �M@      �?              @      B@              @      1@       @     �I@      �?      L@      "@       @              L@     �T@      @      @     �Y@      5@     �d@      D@     @_@     �T@       @              @      ;@      �?              1@      @     �O@      @      E@      2@                      I@     �K@      @      @     �U@      0@     @Y@     �B@     �T@      P@       @              5@      L@      @      "@     �A@      @      c@      4@     �Z@     �A@      �?              @      8@              @      @             �T@      &@      K@      @                       @      ,@              @      �?              3@      "@      @      @                      @      $@                      @             �O@       @      H@      @                      .@      @@      @      @      =@      @     �Q@      "@      J@      =@      �?              "@      2@               @      3@      @     �O@      @      F@      :@                      @      ,@      @      @      $@      �?       @      @       @      @      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���bhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�ܩ���@�	           ��@       	                    �?�Pk�K�@�           �@                          �6@��\)o@�           ��@                            �?0#5e�@�            0z@������������������������       �����O@�            �m@������������������������       ��:ɟ�@o            �f@                            �?P{-s�@�             n@������������������������       �$i��Yq@Y            �`@������������������������       �8+U�	�@F            �Z@
                          �4@CiJ��e	@�           t�@                           @�-(�L@�           (�@������������������������       ���� �@v           ��@������������������������       ��K?4��@             5@                          �9@6�r���	@b           ��@������������������������       �R�z�~t	@j           ؂@������������������������       �L�2��	@�            �y@                            @q�}��E@           `�@                            �?�(��[L@m           `�@                           �?�@���@�             w@������������������������       ���@��?N            �_@������������������������       �N����@�             n@                          �7@�)8�B�@�           @�@������������������������       �,|�|�@�           Ї@������������������������       ��W�xL@�            �m@                           �?��YH@�             p@                           @	'�c@�@V            @a@������������������������       ��Nu"@J             ]@������������������������       �%X	�/@             6@                           @w���6@O            �]@������������������������       �� �rgH @"            �J@������������������������       �M}H*��@-            @P@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     �q@     �@      <@      J@      ~@     �X@     @�@      o@     ؉@     �v@      @@      0@     @h@     @t@      4@     �F@     pv@     �S@     `w@      j@     �y@     @m@      <@              H@     @X@      �?      @     �P@      (@     �d@      I@      d@     �H@      @              9@     �O@               @      ;@      @     �_@     �C@     �Z@      9@      �?               @      A@               @      $@      �?     �Q@      8@      R@      ,@      �?              1@      =@                      1@      @     �K@      .@      A@      &@                      7@      A@      �?      @     �C@      @      D@      &@      K@      8@      @              $@      5@               @      ,@      @      2@      @     �A@      4@      @              *@      *@      �?      @      9@      @      6@      @      3@      @              0@     @b@     `l@      3@      C@     Pr@     �P@      j@     �c@      o@      g@      8@      @     �E@     �P@      @      @      ]@      1@     �[@     �L@      ^@      O@      @      @      C@      P@      @      @      \@      1@      [@     �L@     �]@     �N@       @              @       @                      @               @               @      �?      @      "@     �Y@      d@      ,@     �A@      f@      I@     �X@     @Y@      `@     �^@      1@      @      O@     @X@      "@      :@     �^@      6@      M@     �G@     �T@      O@      (@      @     �D@      P@      @      "@     �K@      <@      D@      K@     �F@     �N@      @             �V@     �k@       @      @     @^@      4@     ��@     �D@     0z@     ``@      @             �T@     �i@      @      @     �Z@      0@     �}@     �A@     pt@     �Z@      @              5@      C@       @              <@      @     �d@       @     �R@      9@                              (@       @              (@      @     �R@      �?      3@      @                      5@      :@                      0@      @     �V@      @      L@      5@                      O@     �d@       @      @     �S@      $@     �s@      ;@     �o@     �T@      @             �B@     @`@       @      @     �I@       @     �p@      1@     �g@      L@      �?              9@      B@               @      <@       @     �E@      $@      P@      :@       @              @      1@      @       @      ,@      @     @U@      @      W@      8@      �?              @      &@       @       @      @       @      G@      �?      I@      .@      �?              @      $@               @      @              D@      �?      G@      "@                              �?       @                       @      @              @      @      �?              @      @       @              "@       @     �C@      @      E@      "@                      �?      �?                      �?       @      9@      @      0@       @                      @      @       @               @              ,@              :@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ>��RhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @3e���f@�	           ��@       	                    �?zE_ �@}           t�@                          �8@��B ��@           ��@                           @
�"dk@{           @�@������������������������       ����k�@            z@������������������������       �v�dx@z            �h@                            @|GL�r�	@�            �m@������������������������       ���.��@Z             a@������������������������       ��]I�
@C             Y@
                           �?V��6k�@e           ��@                           �?���[M	@�           H�@������������������������       ������@�            �p@������������������������       ��Y��	@�           8�@                           �?K����@�            @u@������������������������       ��ٕw(e @8            �V@������������������������       �.��5��@�             o@                           @L�,�Q@.           <�@                          �7@�'��K@�           ��@                           @��j93@>           `�@������������������������       �@�%]�@�            0p@������������������������       �����/� @�           H�@                           @��w�d@�            �o@������������������������       �5M��x�@v            �h@������������������������       ����w��@!            �K@                          �5@v����@Y           (�@                          �1@-'���@�            �r@������������������������       �h2<�@7            �T@������������������������       ��Sf3G$@�             k@                            �?;#�:|@�             o@������������������������       ���`�k@U            @`@������������������������       ��UU���@J            �]@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      r@     ��@     �B@     �M@      {@     @R@      �@     @l@     ȉ@     v@     �A@      6@     `k@     v@      =@      E@     �q@      J@     pw@     �f@      z@     �m@      ;@      "@      Q@      c@      1@      .@     �]@      3@      b@     @P@     �a@      V@      (@       @     �I@      \@      $@      &@      V@       @     @_@     �B@     @\@     �H@      $@      �?     �@@     �M@      $@      @      R@      @     @Z@      .@      U@      :@      �?      �?      2@     �J@              @      0@       @      4@      6@      =@      7@      "@      @      1@     �D@      @      @      >@      &@      4@      <@      >@     �C@       @       @      $@      6@       @              0@      @      *@      5@      .@      =@              @      @      3@      @      @      ,@      @      @      @      .@      $@       @      *@     �b@      i@      (@      ;@     @d@     �@@     �l@     @]@     q@     �b@      .@      *@     �_@     `a@      "@      4@     �`@      8@     �b@      X@     `h@     �^@      ,@              ?@     �D@              @      ?@              K@      "@     �Q@      8@       @      *@     �W@     �X@      "@      0@      Z@      8@     �W@     �U@      _@     �X@      (@              9@     �N@      @      @      ;@      "@     @T@      5@     �S@      ;@      �?              @      @                      @              @@      �?     �C@      @      �?              4@      L@      @      @      8@      "@     �H@      4@     �C@      6@              �?     �Q@     `j@       @      1@      c@      5@     h�@      F@     �y@      ]@       @      �?     �G@     ``@       @      @     �Y@      &@     0|@      5@     �q@     @Q@      @              B@     @Y@       @      @     �O@      &@     �x@      "@     �j@     �D@      @              (@      B@       @              ,@      &@     @[@      @      G@      7@      @              8@     @P@              @     �H@             �q@      @      e@      2@              �?      &@      >@              �?     �C@             �M@      (@     �Q@      <@      @      �?      "@      2@              �?      <@              F@      (@      L@      ;@      @               @      (@                      &@              .@              ,@      �?                      8@      T@      @      (@      I@      $@     @e@      7@     @_@     �G@       @              *@     �C@      �?       @      6@       @     �^@      @      Q@      2@       @              �?      .@              @      @              >@      �?      3@      @       @              (@      8@      �?      @      .@       @     @W@      @     �H@      .@                      &@     �D@      @      @      <@       @     �G@      3@     �L@      =@                      @      ,@                      &@       @      =@      $@      >@      5@                      @      ;@      @      @      1@              2@      "@      ;@       @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��shG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?$0���0@�	           ��@       	                    �?��z-��@           ��@                            �?���I�)@�           H�@                           �?��̎�~@_             d@������������������������       �U+@              J@������������������������       �W`�����??            @[@                           @l�����@-           �~@������������������������       �o�@�            @l@������������������������       �$�M�u@�            `p@
                            �?X�M¸@u           ��@                           @a��Y�9@�            @u@������������������������       ��k�l~0@|             k@������������������������       �o*R�m�@O             _@                          �:@�CLo�@�            �p@������������������������       �\�x��@�             l@������������������������       �$uX��i@            �C@                          �5@�6L�@�           Ȥ@                          �4@!�MK��@�           p�@                           @ls�;YF@�           <�@������������������������       �nqeek@l           ؁@������������������������       ���&�@r           ��@                           �?K�F���@�            �p@������������������������       �Y&Ϩz@F            @Z@������������������������       ���5��@d            �d@                            �?~�^�|I	@            �@                           �?Jt�.�	@�            �u@������������������������       �$<�wQ@O            �_@������������������������       ��'@-�;	@�            �k@                           @gEpT�7	@4           X�@������������������������       ��J���	@n           H�@������������������������       ��9�>xQ@�             r@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        0@     @s@     �@      <@      L@     �y@     @R@     L�@     @l@     ��@      x@      =@             @T@     `e@      @      $@     �X@      &@     �{@     �J@     pr@      T@      @             �B@     �U@       @      @     �F@      @     pp@      A@      _@      F@                      @      6@              �?      (@             @R@      @      C@      @                      @      (@                      @              2@      @      @      @                              $@              �?      @             �K@             �@@      @                      ?@     @P@       @      @     �@@      @     �g@      ?@     �U@      C@                      5@      :@       @      @      7@       @     �M@      9@      B@      =@                      $@     �C@              @      $@      @     ``@      @      I@      "@                      F@      U@      @      @      K@      @     �f@      3@     `e@      B@      @              :@      G@      @       @      ;@      @     �V@      (@     �Z@      3@      @              :@     �@@               @      .@             �B@      &@     �R@      .@      @                      *@      @              (@      @     �J@      �?     �@@      @                      2@      C@              �?      ;@              W@      @      P@      1@                      "@      ?@              �?      1@             �U@      @     �M@      .@                      "@      @                      $@              @      �?      @       @              0@     `l@     �w@      7@      G@     `s@      O@     ��@     �e@     @      s@      :@      @     �U@      k@      @      4@     `a@      8@     �x@      Q@      t@     @b@      $@      @     @R@     �d@      @      &@     @Z@      4@     �u@     �L@     �n@      _@      @      @      G@      V@      @      @     �Q@      0@     �Z@      G@     �Y@     �R@      @              ;@     �S@      �?      @      A@      @     `n@      &@     �a@      I@                      *@      I@      �?      "@      A@      @      G@      &@     �R@      6@      @              @      6@      �?       @      ,@       @      .@      �?      8@      &@      @              "@      <@              �?      4@       @      ?@      $@     �I@      &@      �?      $@     �a@     �c@      2@      :@     `e@      C@     `i@     @Z@      f@      d@      0@             �E@      D@      @      &@     �J@      $@     �P@      D@      B@      D@      @              $@      .@      �?              <@      �?      <@      *@      (@      *@      @             �@@      9@      @      &@      9@      "@      C@      ;@      8@      ;@      �?      $@     �X@     �]@      ,@      .@     �]@      <@      a@     @P@     �a@      ^@      $@      $@     �R@     @U@      ,@      &@     �T@      9@      L@     �M@      R@     �U@      $@              7@      A@              @      B@      @     @T@      @     @Q@      A@        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ��~hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?��tǒr@�	           ��@       	                    @oR@]��@           ��@                           �?�Ӎ���@�           Є@                           �?�p�^&@�            �s@������������������������       ��Õ��@:            �W@������������������������       �laӌ�@�            �k@                          �<@�u���K@�            �u@������������������������       ���S�rb@�            �s@������������������������       � �͓�4@             @@
                           �?�N��%q@u           H�@                           @rS
D1 @�            �u@������������������������       �Z2v�F��?�            `k@������������������������       �nJ��f@N            @_@                          �1@���8Y�@�             n@������������������������       ���>Gtk�?.            @Q@������������������������       �����0@n            �e@                           @MK�,�Y@�           ̤@                          �2@`i�RA�	@�           ��@                           �?گ}�@�            �s@������������������������       �� �'��@             h@������������������������       ����	�p@E             ^@                           �?�mO2�	@           ��@������������������������       ��'h�N@�             t@������������������������       �nV��	
@N           h�@                           @�)9���@�            �@                          �2@�Ke��@�           ��@������������������������       �5��[` @�            �k@������������������������       �G|WE�@g           ��@                           �?Һ��hz@�            �r@������������������������       ���� Q3@S            ``@������������������������       �Ъ�&�@n            `e@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        .@     �s@     p�@     �G@     �O@     �{@     �Q@     ��@     �j@     x�@     �v@     �@@      �?     �V@      f@      @      @      Z@      ,@     {@      H@      r@     �S@      @      �?      R@     �U@       @      @     @S@      "@     �b@      D@     �d@     �L@      @      �?      8@     �C@       @      �?     �G@      @     @S@      ;@      M@      @@      �?      �?      @      "@                      9@              :@      @      3@       @                      5@      >@       @      �?      6@      @     �I@      8@     �C@      8@      �?              H@      H@               @      >@       @     �R@      *@     �Z@      9@       @              E@     �G@              �?      7@       @     @R@       @     �Y@      2@      �?              @      �?              �?      @              �?      @      @      @      �?              2@     �V@       @       @      ;@      @     �q@       @     �_@      5@      @              @      J@               @      0@      @     `f@      @     �Q@      (@                      �?      6@                       @       @     �a@       @     �A@       @                      @      >@               @       @      �?      C@       @     �A@      @                      (@      C@       @              &@       @     �Y@      @      L@      "@      @              @      @                       @              D@      �?      (@              @              "@      ?@       @              "@       @     �O@      @      F@      "@              ,@     �k@     �w@     �E@      M@      u@     �L@     �@     �d@     �~@     �q@      :@      ,@     �e@     �l@     �@@      I@     �m@     �H@     �l@     ``@     �i@      i@      3@      @     �A@     �B@      �?      @      C@             @U@      B@     �C@      A@      �?      @     �@@      1@      �?       @      8@              C@      6@      6@      =@      �?               @      4@              �?      ,@             �G@      ,@      1@      @              $@     �a@      h@      @@     �G@      i@     �H@      b@     �W@     �d@     �d@      2@              $@     �N@      @      2@      K@      @      D@      4@      H@     �J@      @      $@     @`@     �`@      <@      =@     `b@     �E@     @Z@     �R@     @]@     @\@      (@              H@     �b@      $@       @     �X@       @     �u@      B@     r@     @U@      @             �A@      ]@      @      @     �L@      @     �q@      6@     �i@     �I@      @              "@      D@       @              �?      �?     @W@       @      P@       @                      :@      S@       @      @      L@      @     �g@      4@     �a@     �E@      @              *@     �A@      @      @      E@      @      P@      ,@     @U@      A@       @              @      ,@       @       @      5@              7@      @      F@      ,@                      @      5@      @       @      5@      @     �D@      "@     �D@      4@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ���VhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�BX                             �?���{�~@�	           ��@       	                    �?߆L�z�@           8�@                           �?��l��@�           `�@                           �?G�	8��@�            @n@������������������������       �p��4@@             Z@������������������������       ��?g,	@Z            @a@                            @{؄f.�@            �w@������������������������       ���	��]@�            �r@������������������������       ����7̵�?1            �R@
                           �?�a,H@q           �@                            �?�]z��@�            �p@������������������������       �� wZ�@[            `a@������������������������       �ݤܭ3@H            ``@                            �?����
y @�            @u@������������������������       �U�F�9�?<             Z@������������������������       �~��9� @�            �m@                           @Q�
	ei@�           ��@                          �1@9���@�           b�@                           @yQ)�	@�            �t@������������������������       �3�ZPX�@�            �k@������������������������       �_���e@I            �[@                           �?���G�@�           ��@������������������������       �Lt����@           �@������������������������       �v~M?�@�           ��@                           !@�Vũ��	@�            �t@                          �9@q�H��?	@�             s@������������������������       � 92�I	@�            �k@������������������������       ��<3ŀZ@3            �T@������������������������       �H��7zT@             :@�t�bh�h5h8K ��h:��R�(KKKK��h��B�
        =@     Pq@     0�@     �B@     �H@     �{@     �X@     @�@     @k@     ��@     �x@      ;@      �?     �S@     �a@       @      @     �Z@      *@     `{@     �E@     �r@     �V@      @      �?     �B@     �Q@      @      @     �N@      (@     @m@      4@      _@     �H@       @      �?      7@      ?@      @       @      7@      @     �J@      ,@      H@      A@       @      �?      @      &@                      *@              A@      @      :@      $@                      2@      4@      @       @      $@      @      3@      $@      6@      8@       @              ,@      D@              @      C@      @     �f@      @      S@      .@                      "@     �C@              @      @@      @     �a@      @     �J@      *@                      @      �?                      @              C@              7@       @                      E@      R@      @      �?      G@      �?     �i@      7@     �e@     �D@       @             �B@      G@              �?      ?@              J@      0@     �M@      <@                      1@      6@                      "@              8@       @      E@      1@                      4@      8@              �?      6@              <@       @      1@      &@                      @      :@      @              .@      �?      c@      @     �\@      *@       @              �?      @      @              @      �?      K@      �?      @@       @                      @      6@                      $@             �X@      @     �T@      &@       @      <@     �h@     py@      =@     �E@      u@     @U@     ��@     �e@     �~@      s@      7@      0@     �c@      w@      <@      D@     r@     @R@     `@     �a@     �{@     `q@      *@      @      (@      M@              @      :@             @[@      &@     �T@      :@                      "@     �A@              �?      2@             �N@      @     �Q@      4@              @      @      7@               @       @              H@      @      *@      @              *@     @b@     �s@      <@     �B@     pp@     @R@     �x@     ``@     �v@     �o@      *@      @     �D@     `a@      .@      "@     @[@      8@      e@     �E@     �c@     �\@      @      @     @Z@     �e@      *@      <@     @c@     �H@      l@      V@     `i@      a@      @      (@      D@     �B@      �?      @     �G@      (@      N@     �@@     �H@      :@      $@      (@      ?@     �@@      �?      @     �E@      @      N@      @@      H@      9@      "@      @      7@      >@      �?      @      ?@      @     �E@      6@      >@      5@      "@      @       @      @                      (@      @      1@      $@      2@      @                      "@      @                      @      @              �?      �?      �?      �?�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�}-\hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�Bx                             @TTg��E@�	           ��@       	                   �;@�y$I�@d           �@                           �?��2/N@�           Ȝ@                           �?�y��s@p           0�@������������������������       �O��)�8@           p{@������������������������       �8PDG�|@a            �a@                          �3@��I�	@:           ��@������������������������       �ׯ<���@            {@������������������������       �<4��	@,           ��@
                          �A@N��(�	@�            t@                           �?���E��	@�             s@������������������������       ��ɥ1��	@�            0p@������������������������       ��#yP@            �F@������������������������       �(*�ED� @	             1@                           @Gh`@�@6           X�@                           @�тI@�           �@                          �2@��/{A@�           ̒@������������������������       ��IB����?�            �z@������������������������       �:�[`�+@�           H�@������������������������       ���<ܷ@             3@                           @(:�>@C           ��@                           �?�;8�@<           �@������������������������       ��W�D�@}             j@������������������������       �_���\@�             s@������������������������       ��r�u�@             ,@�t�bh�h5h8K ��h:��R�(KKKK��h��B`	        7@     0q@     h�@      C@      H@     p~@     �V@     �@     �h@     �@     `u@      ?@      7@     �j@     `s@      2@      @@     �t@     �P@     �w@     �d@     @v@     �m@      =@       @     �f@      q@      .@      :@     @r@     �H@     �u@     �`@     0t@      e@      6@             �J@      R@       @      @     �S@      @     �e@      4@     ``@     �E@      @              E@      P@       @      @     @P@       @      \@      4@      W@     �@@      @              &@       @                      *@      �?     �N@             �C@      $@               @     �_@      i@      *@      7@     �j@      G@     @f@     �\@      h@     �_@      2@      @      >@     �M@       @      @     �I@      3@      Z@     �B@     �Q@      I@      �?      @     @X@     �a@      &@      1@     `d@      ;@     �R@     �S@     �^@      S@      1@      .@     �@@      C@      @      @      E@      1@      <@      >@     �@@     @Q@      @      "@     �@@     �@@      @      @     �C@      1@      <@      =@     �@@     �P@      @      "@      :@      ;@      @      @      A@      .@      4@      9@      7@     @P@      @              @      @                      @       @       @      @      $@       @      �?      @              @                      @                      �?               @                      O@     �n@      4@      0@      c@      8@     H�@      @@     �{@      Z@       @              E@     �e@      @      @     @W@      0@     `@      0@     Ps@     �O@                      D@     �e@      @      @     @V@      (@     @@      .@     @s@      N@                      &@      N@      @              ,@      �?     �k@      @     @X@      *@                      =@      \@              @     �R@      &@     `q@      &@     `j@     �G@                       @               @              @      @       @      �?      �?      @                      4@     �R@      ,@      *@      N@       @     `b@      0@     �`@     �D@       @              1@     �R@      ,@      "@     �M@      @     `b@      0@      `@     �D@       @              @     �B@      @      @      ,@              T@      @     �F@      $@       @              (@      C@      $@      @     �F@      @     �P@      "@      U@      ?@                      @                      @      �?      @                      @                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ�ohG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                            �5@�)��#*@�	           ��@       	                    @ޗ���j@i           ��@                          �1@�}�:��@`           ��@                           �?N�p{
@�            Pu@������������������������       ��01�@p            �d@������������������������       �݈�i�@w             f@                           @��4�y@y           Ȏ@������������������������       �A��,�@            ��@������������������������       �VlC�X@y            �h@
                          �4@�܀�@	           h�@                           �?2��r�@�           ��@������������������������       �̳��@           �z@������������������������       �Rn���@�            �r@                           @#�w$��@G            @]@������������������������       �~ �u/��?             >@������������������������       ���T�=@2            �U@                           �?t�����@I           8�@                          �<@>�D��V@<           �@                          �9@V�[��p@�            Py@������������������������       ���z� @�            pq@������������������������       �&P�R+�@M            �_@                           @�޿��D@B            �Y@������������������������       �#]�ݼ@/            @S@������������������������       �K��@             :@                           @��c��*	@           H�@                           �?V*�X�
@�           @�@������������������������       �.I[	@�            @j@������������������������       �W;��r%
@z           ��@                           @�s�\�y@           �z@������������������������       �mѷ��%@           py@������������������������       ��N?~�@             3@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        (@     Pp@     ��@      @@     �L@      |@     �X@     �@     �j@     ��@     �w@      8@      @     �X@      s@      ,@      =@     @j@     �C@     P�@     @W@      �@     `b@      @      @     �R@      k@      (@      1@      c@      B@     �v@     @T@     �p@     @X@      @              1@     �O@       @      �?      3@      �?     ``@      5@      L@      >@                      *@      >@       @      �?      ,@      �?      K@      "@      7@      2@                      @     �@@                      @             @S@      (@     �@@      (@              @     �L@      c@      $@      0@     �`@     �A@     �l@      N@     �j@     �P@      @      @      G@     @[@      $@      0@     @]@      8@      f@     �J@      e@      N@      @              &@      F@                      0@      &@      K@      @     �F@      @      @              9@      V@       @      (@      M@      @      v@      (@     `n@      I@                      6@     �O@       @      (@      J@      �?     �s@      "@      j@     �E@                      "@      B@      �?       @      C@      �?      h@      @      Z@      >@                      *@      ;@      �?      @      ,@             �^@      @     @Z@      *@                      @      9@                      @       @     �B@      @      A@      @                      �?       @                      @              ,@              $@                               @      7@                      @       @      7@      @      8@      @              "@     @d@      l@      2@      <@      n@      N@     �s@     �]@     �s@      m@      1@             �F@     �S@              @     �H@      @      ^@      9@     @^@     �K@      @             �D@     @P@              �?      D@      @      Z@      .@     �Y@      =@       @              =@     �@@              �?      ?@       @     �T@      @      Q@      8@       @              (@      @@                      "@      @      6@       @     �A@      @                      @      *@              @      "@      �?      0@      $@      2@      :@       @              @      $@              @      "@              @      "@      "@      7@       @                      @                              �?      "@      �?      "@      @              "@     @]@     @b@      2@      7@     �g@      K@      h@     �W@     �h@     @f@      *@      "@     @W@     @Y@      1@      4@      \@     �H@     �W@     @T@     @W@     �_@      *@              (@      4@      @      "@     �@@      @      ?@      7@      <@      D@       @      "@     @T@     @T@      &@      &@     �S@     �E@     �O@      M@     @P@     �U@      &@              8@     �F@      �?      @     �S@      @     �X@      *@     @Z@      J@                      6@     �E@              @     �Q@      @     @X@      &@      Z@      J@                       @       @      �?               @      �?       @       @      �?                �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ �uIhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @iD^��R@�	           ��@       	                    �?������@n           p�@                           �?�ӹ#�@�           ��@                           �?6���@%            }@������������������������       ������@            `i@������������������������       ���Q��@�            pp@                          �<@'��y�@z            @h@������������������������       �cY�8� @s             g@������������������������       �QcX^@             $@
                           �?Iu����	@�           ��@                          �3@��$�E@           p}@������������������������       �J;O�g@V            �c@������������������������       ����Q@�            �s@                           @����	@�           4�@������������������������       �yZ̦�	@a           Ѝ@������������������������       ��Z��@Y            `b@                          �4@��^��@8           D�@                           �?��C�Ir@K           �@                           �?�=�2�?�            �u@������������������������       ��}EX�?�            �h@������������������������       ��EW�G�?]            @b@                          �1@0��]n@k           X�@������������������������       ���iw�?�             k@������������������������       ����
��@�             w@                            �?g��%@�           p�@                          �5@�&q�R@
           �x@������������������������       �OUD���@;            �V@������������������������       �̎�P@�            �r@                           @И2��@�            Pv@������������������������       �9.W6G	@�             l@������������������������       �	+4Q_@R            �`@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        2@     Ps@     8�@      <@      M@     �|@     �W@     0�@     �i@     Ȉ@     �v@      ?@      0@     �l@     �r@      7@     �F@     @s@     @S@     �y@     �d@      w@     Pp@      :@       @     �L@     �S@              "@     �P@      @     @g@      7@     �d@      P@      �?       @     �D@     @P@               @     �M@      @     @X@      3@     �\@     �J@      �?       @      ,@      4@              @      @@      @      I@       @     �E@      8@                      ;@     �F@              @      ;@             �G@      &@      R@      =@      �?              0@      ,@              �?       @      �?     @V@      @      I@      &@                      0@      (@              �?      @      �?      V@      �?     �H@      &@                               @                      @              �?      @      �?                      ,@     �e@      l@      7@      B@      n@     �Q@     �k@     �a@     �i@     �h@      9@      �?      @@      S@      @      .@     @T@      &@     @V@      =@     �R@     �J@      @      �?      6@      8@                      7@      @     �D@      @      9@      $@      �?              $@      J@      @      .@      M@       @      H@      6@      I@     �E@      @      *@     �a@     �b@      4@      5@      d@     �M@     �`@     @\@     @`@      b@      3@       @      `@     @_@      4@      5@      a@     �K@     �Z@     �T@     �^@     �`@      ,@      @      (@      7@                      7@      @      <@      >@      @      $@      @       @      T@      k@      @      *@      c@      2@     ��@      D@     pz@     �X@      @              >@      [@       @      @      O@      @      {@      1@      m@      D@                      (@      ?@              �?      ,@              i@      @     @P@      .@                      "@      0@              �?      "@             @]@      @      ?@      (@                      @      .@                      @              U@       @      A@      @                      2@     @S@       @      @      H@      @     �l@      (@     �d@      9@                      @      9@              �?      *@              W@      �?     @S@      @                      ,@      J@       @      @     �A@      @     `a@      &@     �V@      5@               @      I@      [@      @       @     �V@      .@     `h@      7@     �g@     �M@      @              9@     @P@              @      F@      &@     �Y@      1@     �V@     �@@      �?                      :@              �?      @      @      ;@      �?      6@       @      �?              9@     �C@              @     �B@      @     �R@      0@     @Q@      ?@               @      9@     �E@      @      @     �G@      @     @W@      @      Y@      :@      @       @      $@      8@              �?      ?@      @     �R@       @     �N@      ,@      �?              .@      3@      @      @      0@      �?      2@      @     �C@      (@      @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJ:��9hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�)Ca1@�	           ��@       	                    �?����&@�           �@                          �6@�><mѳ@t           ��@                            @�D��o@           py@������������������������       �`�ُ͐@�            s@������������������������       �Ƨ,��@C            �Y@                           �?H2�_Jr@i            �d@������������������������       �J�)6�@-            @R@������������������������       �]�o��@<            �W@
                          �2@�x͌:@�           0�@                          �1@�c�� @�            @l@������������������������       ���!�1Z�?Q            @a@������������������������       �3�)� @2             V@                            �?���/�t@           @z@������������������������       ��1�9�@�            �l@������������������������       ��A�/�@x            �g@                          �4@���)1@�           
�@                           @�&	_ �@            ��@                           @�P���@           Ȉ@������������������������       ����;pl@           `y@������������������������       �������@            0x@                           �?v�oc~@�            `y@������������������������       ��5%���@n            �f@������������������������       �$���@�             l@                           @Єr��`	@�           X�@                          �8@��J�a	@:           \�@������������������������       �"G�BR@�           0�@������������������������       �z��E�	@y           ��@                           �?�d;gL�	@�            �g@������������������������       �KG]@             =@������������������������       �a5A�|�	@p            @d@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        9@     `s@     @�@      ?@      I@     z@     @Q@     T�@     �k@     `�@     �u@      @@             �U@     �f@      @       @     �X@      @     p{@      A@     `q@     �U@      @              =@     �S@      @      @      I@      @     �m@      2@      [@     �D@                      *@      N@      �?       @     �A@      @      h@      *@      P@      7@                      @      H@      �?       @      6@      @      c@      &@     �H@      (@                      "@      (@                      *@              D@       @      .@      &@                      0@      2@       @      @      .@              G@      @      F@      2@                      @      $@       @      @      (@              @      @      5@      &@                      &@       @                      @             �D@      �?      7@      @                     �L@     �Y@              @     �H@      �?      i@      0@     @e@     �F@      @              @      :@                      ,@             @[@       @     �N@       @      �?              @      0@                      "@             @S@      �?      <@      @      �?               @      $@                      @              @@      �?     �@@      @                      J@      S@              @     �A@      �?     �V@      ,@     @[@     �B@       @              8@      F@              @      (@      �?     �D@      "@      Q@      9@       @              <@      @@                      7@              I@      @     �D@      (@              9@      l@     @w@      <@      E@     �s@     @P@     ��@     �g@     ��@     `p@      =@      @     �P@     @e@      "@      (@     �[@      $@     Pw@     @Q@     �p@     @Y@      @      @      F@      Z@      @       @     �V@      @     @l@      B@      h@     @S@      �?      @      9@      J@      @      @      O@      @      S@     �@@     @U@     �L@      �?              3@      J@      �?      @      =@       @     �b@      @     �Z@      4@              �?      6@     �P@      @      @      3@      @     `b@     �@@      S@      8@      @              ,@      =@       @      @       @      @     @Q@      .@      2@      2@      �?      �?       @     �B@      �?              &@      �?     �S@      2@      M@      @      @      5@     �c@     @i@      3@      >@      j@     �K@      m@     �]@     �p@      d@      6@      1@      a@     @e@      ,@      =@     �f@     �H@      j@     �V@     �n@     �b@      (@       @      S@     �Z@      @      0@     �[@      6@     @`@      ?@     �`@      Q@      @      "@     �N@     �O@      $@      *@     �Q@      ;@     �S@      N@     @\@     @T@      @      @      5@      @@      @      �?      :@      @      9@      <@      5@      (@      $@              @       @                      $@                       @      �?      @              @      2@      >@      @      �?      0@      @      9@      4@      4@      @      $@�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJlQP;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�\��Xi@�	           ��@       	                   �3@�jߗ<	@�           �@                           @WEt.�@           �|@                           �?���c�|@�             t@������������������������       �����@O            ``@������������������������       ���]dN@s            �g@                           @S�WUA@]             a@������������������������       ����77@K            �[@������������������������       ��bn�@             :@
                          �;@I�E��	@�           Ē@                           �?%Sc�m	@1           ��@������������������������       ���x	@�            �w@������������������������       �&���	@X           ��@                          �<@j��%�Z	@�            �o@������������������������       ���(�@&            @P@������������������������       ���Z%/�@u            �g@                           @�Xi�J$@�           ��@                          �2@�>t��A@|           (�@                          �1@�{���/@�            �p@������������������������       �Mq��� @i            �d@������������������������       �A��
�d@E            �Z@                           @��7"@�           ��@������������������������       �o��%�@           �z@������������������������       ��_��!@�            �r@                           �?�����@-           ��@                            @�'��Z�@           0{@������������������������       �ۍ�2�c@�            0w@������������������������       ��y]�*�?,             P@                           @dV@��@           ��@������������������������       ��]C �@�           0�@������������������������       �dz��@E            @\@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        6@     Pr@     �@      ;@      N@     0{@     �S@     h�@     �i@     ��@     �y@     �@@      4@      f@     @p@      3@      A@     �m@     �F@     `m@     �]@      p@     �l@      =@      @      >@      Q@       @       @      Q@      @      \@      6@     �T@     �L@      @      �?      &@      H@      �?       @      E@      @     �U@      *@     �Q@      E@              �?      �?      4@      �?              6@      �?      D@       @      8@      *@                      $@      <@               @      4@       @     �G@      @      G@      =@              @      3@      4@      �?              :@      �?      9@      "@      *@      .@      @       @      3@      1@      �?              3@              7@      "@      &@      "@      �?      �?              @                      @      �?       @               @      @      @      0@     `b@      h@      1@      @@      e@     �D@     �^@      X@     �e@     `e@      8@      @     �\@     �b@      .@      9@     �a@      <@     �Z@     �R@      c@     �[@      5@              N@     �P@      $@       @     �G@      0@      B@      @@      G@      H@      "@      @      K@      U@      @      1@     �W@      (@     �Q@     �E@     �Z@     �O@      (@      &@     �@@     �D@       @      @      <@      *@      0@      5@      4@      N@      @      "@      "@      @       @              @      @      $@              @      &@      �?       @      8@      A@              @      5@      "@      @      5@      .@     �H@       @       @      ]@     �s@       @      :@     �h@     �@@     �@     �U@     ��@      g@      @       @      N@     @d@       @      "@      \@      :@     Pq@      L@      j@     @T@      �?              @      G@              �?      4@             �]@      *@      H@      5@                       @      5@                      $@             �T@      *@      =@      @                      �?      9@              �?      $@              B@              3@      ,@               @     �L@      ]@       @       @      W@      :@     �c@     �E@      d@      N@      �?       @      ;@      K@              @      P@      2@      \@      1@      W@      C@      �?              >@      O@       @      @      <@       @      G@      :@     @Q@      6@                      L@     �c@      @      1@     �U@      @     �|@      ?@     �t@      Z@      @               @      I@              @      5@       @     @i@      $@     �Z@      >@      �?               @     �H@              @      4@       @     �c@       @     �V@      >@      �?                      �?              �?      �?             �E@       @      0@                              H@     �Z@      @      (@     @P@      @     0p@      5@      l@     �R@       @              E@     �W@      @      (@      K@      @     �k@      ,@     �h@      P@                      @      (@      �?              &@             �B@      @      ;@      $@       @�t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJi>DhG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             @�����8@�	           ��@       	                     @Yu��D�@�           <�@                            �?\�r�@l           ��@                           �?�7[sB�@�           �@������������������������       ���8�d{@            z@������������������������       �ƠK6R�@�           (�@                           �?�ǐ3��@�            �k@������������������������       ���+L�@.             Q@������������������������       ���8�9}@[            `c@
                           �?W�y���@           ��@                           �?C��@�            �j@������������������������       ��״�̱@D            �Z@������������������������       ���wx��@R            �Z@                           �?�?ROk	@�           �@������������������������       ��?d��q	@�            �j@������������������������       �zX,G�@�            �x@                          �7@�c�k�@B           ��@                           �?�eW�~@>           $�@                           @Ȼ��:�?+           �~@������������������������       ���^�?�            �t@������������������������       ������@^             c@                          �1@|׽���@           �@������������������������       �>�Cu� @{            �g@������������������������       �n�W�@�           �@                            @#�n�@            z@                           @���
@�            �t@������������������������       �Q���W�@�            �j@������������������������       �{a�x�@J             ^@                           �??���@2            �U@������������������������       �g���j��?             D@������������������������       �\%����@             G@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        7@      s@     ��@      :@     �N@     }@     �T@     �@     `h@     P�@      w@      8@      6@      l@     �s@      1@     �I@     �t@     @Q@      x@     �d@     pv@      o@      3@       @     �`@     �g@      &@      ?@     @j@     �I@     �m@     �\@     @n@     @b@      $@       @      ]@      d@      &@      =@     �c@      D@      i@     @X@     `j@     �]@      "@      �?      A@     @Q@      @      @     �L@      ,@     �Q@     �E@      Q@      H@      @      @     �T@      W@       @      7@     �Y@      :@      `@      K@     �a@     �Q@      @              0@      =@               @     �I@      &@      B@      2@      ?@      <@      �?              @      @                      &@      @      ,@      @      &@      $@                      &@      6@               @      D@       @      6@      &@      4@      2@      �?      ,@      W@     �^@      @      4@     @^@      2@     �b@      J@     @]@     �Y@      "@              7@      A@      �?      @      6@       @     �P@       @      A@      2@                      $@      .@      �?      @      $@       @     �C@       @      0@       @                      *@      3@              �?      (@              ;@      @      2@      $@              ,@     @Q@     @V@      @      .@     �X@      0@      U@      F@     �T@      U@      "@      @      ;@     �A@      @      "@      A@      @      =@      @      7@      A@      @      "@      E@      K@      �?      @     @P@      $@     �K@      D@      N@      I@      @      �?      T@     �j@      "@      $@     �`@      ,@      �@      <@     0|@      ^@      @             �J@      e@      @      @     �V@      (@     ��@      &@     �t@     �Q@      @              *@      L@              �?      6@       @     0p@       @     �\@      2@      �?               @     �A@                      $@       @     �g@              T@      $@                      @      5@              �?      (@             @Q@       @      A@       @      �?              D@     @\@      @      @      Q@      $@     Pq@      "@     `k@     �J@       @              �?      9@              �?      ,@              T@              N@      $@                     �C@      V@      @      @      K@      $@     �h@      "@     �c@     �E@       @      �?      ;@      G@      @      @      F@       @      Z@      1@     �]@     �H@       @      �?      :@      E@       @      @      C@       @     �N@      &@     �Y@      E@       @      �?      ,@      >@              @      8@              F@      @      O@      ;@       @              (@      (@       @              ,@       @      1@      @      D@      .@                      �?      @       @      �?      @             �E@      @      0@      @                      �?                                              9@      @      @      @                              @       @      �?      @              2@      �?      $@      @        �t�bubhhubh)��}�(hh.hhhKhKhKhG        hhMhNhJϛ;hG        hNhG        h0Kh1Kh2h5h8K ��h:��R�(KK��hT�C`              �?       @      @      @      @      @      @       @      "@      $@      &@�t�bhGhYh\C       ���R�haKhbheKh5h8K ��h:��R�(KK��h\�C       �t�bK��R�}�(hKhoKhph5h8K ��h:��R�(KK��hw�B�                             �?�{dt}@�	           ��@       	                    �?�����@�           Ԓ@                           �?���#{3@'           }@                            �?/|��Y:@�            `h@������������������������       ��\�<:@Q            @_@������������������������       ��ik@/            �Q@                            �?Gݾ.#�@�            �p@������������������������       ������@1            �S@������������������������       �G���#@v            �g@
                           �?ܧ�s�@�            �@                            �?K�Te�N@           `{@������������������������       �YHSޭ�@<            �V@������������������������       �8w���@�            �u@                          �4@,��ͽ@�            �r@������������������������       �6'X�� @y            �g@������������������������       �ُ�1�@H             \@                          �3@�Hes�C@�           (�@                          �1@���D6�@E           ��@                           @A+g!��@�            �w@������������������������       ��!� �6@%            �I@������������������������       ��}�8�@�            �t@                            @W���
@T           ��@������������������������       �Ԉ�!�L@�             x@������������������������       ����hĶ@d            �b@                           @���	@n           �@                            �?��ep�	@�           `�@������������������������       �%L�Ts	@�            `s@������������������������       ������	@            �@                           @��8vj9@�           X�@������������������������       �<楢�@!           �|@������������������������       �S>��e�@�             l@�t�bh�h5h8K ��h:��R�(KKKK��h��B�        4@     `r@     p�@      B@     �L@      {@      T@     �@     �o@     P�@     Pu@      C@       @     �T@     �d@              2@      X@      ,@     py@     �G@     `r@     @Q@      "@       @      K@      S@              ,@     �H@      �?     �W@      <@     �Y@      D@      @       @      0@      9@                      6@             �J@      "@     �J@      *@       @       @      "@      1@                      0@              A@       @      @@      &@       @              @       @                      @              3@      @      5@       @                      C@     �I@              ,@      ;@      �?     �D@      3@     �H@      ;@      @              @      2@              @      $@              .@      @      4@      @                     �@@     �@@              &@      1@      �?      :@      .@      =@      7@      @              <@     �V@              @     �G@      *@     �s@      3@      h@      =@      @              0@      K@              @      >@      @     �i@      (@     @W@      2@                              *@              @      @      @      F@              0@      @                      0@     �D@              �?      8@      �?      d@      (@     @S@      .@                      (@     �B@                      1@      @     @[@      @     �X@      &@      @              $@      7@                      @             �U@      �?     �J@      @      @               @      ,@                      $@      @      6@      @      G@      @      �?      2@     �j@     px@      B@     �C@      u@     �P@     `�@     �i@      �@      q@      =@      @     �D@     @^@       @      "@     �T@      &@      q@     �I@     �k@     @V@      @              ,@      K@      @      @      ;@             �a@      (@     �W@      >@                      @       @                       @              5@      @      @      @                      "@      J@      @      @      9@             @^@      @     �U@      7@              @      ;@     �P@      @      @      L@      &@     @`@     �C@      `@     �M@      @              4@     �I@      @       @      @@      @     �Z@      <@     �W@     �B@      @      @      @      0@              @      8@      @      8@      &@      A@      6@              .@     `e@     �p@      <@      >@     �o@     �K@     �s@     @c@     `r@     �f@      :@      *@      ^@     �e@      5@      7@     `h@     �F@     �Z@     �^@     `b@     @^@      7@              F@      C@      @      "@      N@      ,@      E@      C@      :@      9@      @      *@      S@      a@      ,@      ,@     �`@      ?@      P@     @U@     @^@      X@      0@       @     �I@     �W@      @      @      M@      $@     @j@      ?@     `b@      O@      @       @      ?@     �N@              @      D@      @     �c@      ,@     @Z@      B@      @              4@      A@      @      @      2@      @      J@      1@      E@      :@        �t�bubhhubehhub.