��R0      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K �min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�CP                                                                	       �t�b�
n_classes_�h�scalar���h%C
       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h%�C
       �t�bK��R�}�(h	K
�
node_count�KS�nodes�hhK ��h��R�(KKS��h"�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hHh%K ��hIh%K��hJh%K��hKh"�f8�����R�(Kh&NNNJ����J����K t�bK��hLhVK ��hMh%K(��hNhVK0��uK8KKt�b�B(         :                   �7@�p.0�w�?�             e@                           �?B���?t             ]@                           @�m��?��?&             C@                          �4@h/�����?             ;@                          �3@k��\��?             1@                            �?p=
ףp�?
             $@������������������������       �                     @       	                    �?�8��8��?             @������������������������       �                     @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �      �?              @                           �?0�����?             @������������������������       �      �?              @������������������������       �                     @                          �6@��(\���?
             $@                          �5@�����H�?	             "@������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           �?F]t�E�?             &@������������������������       �                     @                          �6@:/����?             @                           @{�G�z�?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @        3                     @w��"�?N            �S@!       2                     �?#��Q��??            �O@"       -                    @VUUUUU�?$             B@#       ,                    @
ףp=
�?             4@$       %                     �?&�q-�?             *@������������������������       �                     �?&       +                    �?      �?             (@'       *                   �2@���Q��?
             $@(       )                    �?X�<ݚ�?	             "@������������������������       �      �?             @������������������������       ����Q��?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @.       /                    @     ��?             0@������������������������       �                     *@0       1                    !@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@4       7                    @6�h$��?             .@5       6                   �1@�q�q�?             @������������������������       �                      @������������������������       �                     �?8       9                   �5@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?;       P                     @�9J����?4             J@<       K                    :@ʤ��IF�?!            �@@=       D                     �?:/����?             ,@>       ?                    �?0�����?             @������������������������       �                     @@       A                    @VUUUUU�?             @������������������������       �                     �?B       C                   �8@      �?              @������������������������       �                     �?������������������������       �                     �?E       J                   �8@�$I�$I�?             @F       G                    @�q�q�?             @������������������������       �                      @H       I                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?L       O                   �<@�S����?             3@M       N                     �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@Q       R                    �?�KM�]�?             3@������������������������       �                      @������������������������       �                     1@�t�b�values�hhK ��h��R�(KKSKK
��hV�B�        *@      G@      ?@       @      1@      4@       @      >@      �?      @      (@      E@      6@       @                       @      >@              @      $@              .@       @                       @      @              @       @              .@                               @       @                      @              @                               @      �?                       @              @                              �?                                              @                                                               @              @                              �?                                              @                                                               @                                              �?                              �?                                                                              �?                                              �?                              @                                              �?      �?                                                                      �?      �?                      @                                                                              �?               @                                      �?                      �?               @                                                                              @                                                              �?              �?                                                                              �?                                                              �?                                                                                                                                      �?                       @                       @                              @              @                                                                              @       @                       @                              @                       @                       @                              �?                       @                                                      �?                                                                              �?                       @                                                                                                       @                                                                                                               @                       @      E@      @                                      9@               @             �D@      @                                      ,@               @              ,@      @                                      ,@               @              �?      @                                      *@                              �?      @                                      @                              �?                                                                                      @                                      @                                      @                                      @                                      @                                      @                                       @                                       @                                      @                                       @                                      �?                                                                                                                       @                                                                              @                              *@                                              �?               @              *@                                                                                                                              �?               @                                                              �?                                                                                               @              ;@                                                                       @      �?      �?                                      &@                       @      �?                                                                       @                                                                                      �?                                                                                      �?                                      &@                                                                              &@                                      �?                                                              �?      @      "@              1@      4@                      �?              �?      @      @              1@      @                      �?              �?      @      @              �?                              �?              �?              @                                              �?                              @                                                              �?              �?                                              �?                                                                              �?              �?              �?                                                              �?                                                                                              �?                                                                      @       @              �?                                                      @       @                                                                       @                                                                               @       @                                                                       @                                                                                       @                                                                                              �?                                                                              0@      @                                                                       @      @                                                                              @                                                                       @                                                                              ,@                                                               @                      1@                                                       @                                                                                                      1@                                �t�bub�_sklearn_version��1.1.0�ub.